magic
tech sky130A
magscale 1 2
timestamp 1685633567
<< metal1 >>
rect 62 2368 3546 2378
rect 3636 2368 4024 2400
rect 62 2340 4024 2368
rect 62 2308 3696 2340
rect 62 2306 3546 2308
rect -514 2200 3310 2260
rect -514 132 -454 2200
rect -218 2052 3562 2132
rect -218 1402 -128 2052
rect 3472 1402 3562 2052
rect -218 1270 3562 1402
rect -214 940 3566 1066
rect -214 290 -122 940
rect 3478 290 3566 940
rect -214 204 3566 290
rect -514 130 154 132
rect -514 72 3312 130
rect 86 70 3312 72
rect 58 26 3616 28
rect 58 -26 104 26
rect 3288 22 3616 26
rect 3964 22 4024 2340
rect 3288 -26 4024 22
rect 58 -38 4024 -26
<< via1 >>
rect -128 1402 3472 2052
rect -122 290 3478 940
rect 104 -26 3288 26
<< metal2 >>
rect -192 2756 3540 2894
rect -192 2194 -18 2756
rect 3332 2392 3540 2756
rect 3322 2304 3532 2392
rect 3332 2198 3540 2304
rect 3322 2194 3540 2198
rect -192 2132 3540 2194
rect -218 2052 3562 2132
rect -218 1402 -128 2052
rect 3472 1402 3562 2052
rect -218 1270 3562 1402
rect -214 940 3566 1066
rect -214 290 -122 940
rect 3478 290 3566 940
rect -214 234 3566 290
rect -214 204 -36 234
rect -206 -324 -36 204
rect 3300 204 3566 234
rect 3300 -264 3536 204
rect 3300 -324 3526 -264
rect -206 -394 3526 -324
<< via2 >>
rect -18 2392 3332 2756
rect -18 2304 3322 2392
rect -18 2198 3332 2304
rect -18 2194 3322 2198
rect -36 26 3300 234
rect -36 -26 104 26
rect 104 -26 3288 26
rect 3288 -26 3300 26
rect -36 -324 3300 -26
<< metal3 >>
rect -204 2756 3526 2892
rect -204 2742 -18 2756
rect -204 2204 -26 2742
rect 3332 2392 3526 2756
rect 3322 2304 3526 2392
rect -204 2194 -18 2204
rect 3332 2198 3526 2304
rect 3322 2194 3526 2198
rect -204 2040 3526 2194
rect -204 234 3526 272
rect -204 -324 -36 234
rect 3300 -324 3526 234
rect -204 -580 3526 -324
<< via3 >>
rect -26 2204 -18 2742
rect -18 2204 3310 2742
rect 4 -324 3288 170
<< metal4 >>
rect 4712 3236 6226 3258
rect -2424 186 -1112 3172
rect -512 2742 6226 3236
rect -512 2204 -26 2742
rect 3310 2204 6226 2742
rect -512 2000 6226 2204
rect 4348 1890 6226 2000
rect 4712 1770 6226 1890
rect -418 186 4348 220
rect -2424 170 4348 186
rect -2424 -324 4 170
rect 3288 -324 4348 170
rect -2424 -1232 4348 -324
rect -2424 -1256 -36 -1232
rect -2424 -1262 -1112 -1256
use sky130_fd_pr__pfet_01v8_7HKEJJ  sky130_fd_pr__pfet_01v8_7HKEJJ_0
timestamp 1684691938
transform 1 0 1694 0 1 1166
box -1747 -1219 1747 1219
<< end >>
