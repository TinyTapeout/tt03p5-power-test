VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_power_test
  CLASS BLOCK ;
  FOREIGN tt_um_power_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 107.800 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 107.800 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 107.260 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 105.220 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 107.260 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 105.220 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 107.260 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 105.220 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 107.260 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 107.800 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 107.260 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 107.260 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 102.500 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 107.260 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 107.260 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 104.540 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 107.260 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 107.800 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 100.460 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 102.500 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 104.540 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 102.500 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 102.500 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 102.500 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 102.500 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 100.460 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 101.820 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 107.260 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 107.260 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 100.460 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 107.260 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 107.260 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 100.460 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 100.460 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 107.260 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 107.260 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 106.580 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 107.260 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 107.260 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 107.260 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 106.580 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 107.260 66.850 108.800 ;
    END
  END uo_out[7]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.930 5.200 45.530 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.140 5.200 84.740 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.350 5.200 123.950 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 161.560 5.200 163.160 103.600 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.250 -2.010 2.775 103.130 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 6.225 -13.250 8.325 -3.150 ;
      LAYER nwell ;
        RECT 8.345 -13.295 69.175 -3.115 ;
      LAYER li1 ;
        RECT 5.520 0.000 162.380 103.445 ;
        RECT 8.680 -3.295 68.840 -3.290 ;
        RECT 6.405 -3.500 8.145 -3.330 ;
        RECT 6.405 -4.190 6.575 -3.500 ;
        RECT 7.055 -4.010 7.485 -3.840 ;
        RECT 6.955 -4.190 7.125 -4.180 ;
        RECT 6.405 -9.110 7.125 -4.190 ;
        RECT 6.400 -11.250 7.125 -9.110 ;
        RECT 6.405 -12.220 7.125 -11.250 ;
        RECT 7.425 -12.220 7.595 -4.180 ;
        RECT 6.405 -12.900 6.575 -12.220 ;
        RECT 7.115 -12.560 7.455 -12.390 ;
        RECT 7.975 -12.900 8.145 -3.500 ;
        RECT 6.405 -13.070 8.145 -12.900 ;
        RECT 8.525 -3.470 68.995 -3.295 ;
        RECT 8.525 -12.945 8.695 -3.470 ;
        RECT 9.185 -3.955 9.565 -3.755 ;
        RECT 10.095 -4.180 10.265 -3.470 ;
        RECT 11.305 -3.965 11.635 -3.795 ;
        RECT 12.265 -3.965 12.595 -3.795 ;
        RECT 13.225 -3.965 13.555 -3.795 ;
        RECT 14.185 -3.965 14.515 -3.795 ;
        RECT 15.145 -3.965 15.475 -3.795 ;
        RECT 16.105 -3.965 16.435 -3.795 ;
        RECT 17.065 -3.965 17.395 -3.795 ;
        RECT 18.025 -3.965 18.355 -3.795 ;
        RECT 18.985 -3.965 19.315 -3.795 ;
        RECT 19.945 -3.965 20.275 -3.795 ;
        RECT 20.905 -3.965 21.235 -3.795 ;
        RECT 21.865 -3.965 22.195 -3.795 ;
        RECT 22.825 -3.965 23.155 -3.795 ;
        RECT 23.785 -3.965 24.115 -3.795 ;
        RECT 24.745 -3.965 25.075 -3.795 ;
        RECT 25.705 -3.965 26.035 -3.795 ;
        RECT 26.665 -3.965 26.995 -3.795 ;
        RECT 27.625 -3.965 27.955 -3.795 ;
        RECT 28.585 -3.965 28.915 -3.795 ;
        RECT 29.545 -3.965 29.875 -3.795 ;
        RECT 30.505 -3.965 30.835 -3.795 ;
        RECT 31.465 -3.965 31.795 -3.795 ;
        RECT 32.425 -3.965 32.755 -3.795 ;
        RECT 33.385 -3.965 33.715 -3.795 ;
        RECT 34.345 -3.965 34.675 -3.795 ;
        RECT 35.305 -3.965 35.635 -3.795 ;
        RECT 36.265 -3.965 36.595 -3.795 ;
        RECT 37.225 -3.965 37.555 -3.795 ;
        RECT 38.185 -3.965 38.515 -3.795 ;
        RECT 39.145 -3.965 39.475 -3.795 ;
        RECT 40.095 -3.965 40.425 -3.795 ;
        RECT 41.055 -3.965 41.385 -3.795 ;
        RECT 42.015 -3.965 42.345 -3.795 ;
        RECT 42.975 -3.965 43.305 -3.795 ;
        RECT 43.935 -3.965 44.265 -3.795 ;
        RECT 44.895 -3.965 45.225 -3.795 ;
        RECT 45.855 -3.965 46.185 -3.795 ;
        RECT 46.815 -3.965 47.145 -3.795 ;
        RECT 47.775 -3.965 48.105 -3.795 ;
        RECT 48.735 -3.965 49.065 -3.795 ;
        RECT 49.695 -3.965 50.025 -3.795 ;
        RECT 50.655 -3.965 50.985 -3.795 ;
        RECT 51.615 -3.965 51.945 -3.795 ;
        RECT 52.575 -3.965 52.905 -3.795 ;
        RECT 53.535 -3.965 53.865 -3.795 ;
        RECT 54.495 -3.965 54.825 -3.795 ;
        RECT 55.455 -3.965 55.785 -3.795 ;
        RECT 56.415 -3.965 56.745 -3.795 ;
        RECT 57.375 -3.965 57.705 -3.795 ;
        RECT 58.335 -3.965 58.665 -3.795 ;
        RECT 59.295 -3.965 59.625 -3.795 ;
        RECT 60.255 -3.965 60.585 -3.795 ;
        RECT 61.215 -3.965 61.545 -3.795 ;
        RECT 62.175 -3.965 62.505 -3.795 ;
        RECT 63.135 -3.965 63.465 -3.795 ;
        RECT 64.095 -3.965 64.425 -3.795 ;
        RECT 65.055 -3.965 65.385 -3.795 ;
        RECT 66.015 -3.965 66.345 -3.795 ;
        RECT 66.975 -3.965 67.305 -3.795 ;
        RECT 67.935 -3.965 68.265 -3.795 ;
        RECT 9.570 -4.185 10.265 -4.180 ;
        RECT 9.095 -12.225 9.265 -4.185 ;
        RECT 9.535 -12.225 10.265 -4.185 ;
        RECT 10.665 -12.225 10.835 -4.185 ;
        RECT 11.145 -12.225 11.315 -4.185 ;
        RECT 11.625 -12.225 11.795 -4.185 ;
        RECT 12.105 -12.225 12.275 -4.185 ;
        RECT 12.585 -12.225 12.755 -4.185 ;
        RECT 13.065 -12.225 13.235 -4.185 ;
        RECT 13.545 -12.225 13.715 -4.185 ;
        RECT 14.025 -12.225 14.195 -4.185 ;
        RECT 14.505 -12.225 14.675 -4.185 ;
        RECT 14.985 -12.225 15.155 -4.185 ;
        RECT 15.465 -12.225 15.635 -4.185 ;
        RECT 15.945 -12.225 16.115 -4.185 ;
        RECT 16.425 -12.225 16.595 -4.185 ;
        RECT 16.905 -12.225 17.075 -4.185 ;
        RECT 17.385 -12.225 17.555 -4.185 ;
        RECT 17.865 -12.225 18.035 -4.185 ;
        RECT 18.345 -12.225 18.515 -4.185 ;
        RECT 18.825 -12.225 18.995 -4.185 ;
        RECT 19.305 -12.225 19.475 -4.185 ;
        RECT 19.785 -12.225 19.955 -4.185 ;
        RECT 20.265 -12.225 20.435 -4.185 ;
        RECT 20.745 -12.225 20.915 -4.185 ;
        RECT 21.225 -12.225 21.395 -4.185 ;
        RECT 21.705 -12.225 21.875 -4.185 ;
        RECT 22.185 -12.225 22.355 -4.185 ;
        RECT 22.665 -12.225 22.835 -4.185 ;
        RECT 23.145 -12.225 23.315 -4.185 ;
        RECT 23.625 -12.225 23.795 -4.185 ;
        RECT 24.105 -12.225 24.275 -4.185 ;
        RECT 24.585 -12.225 24.755 -4.185 ;
        RECT 25.065 -12.225 25.235 -4.185 ;
        RECT 25.545 -12.225 25.715 -4.185 ;
        RECT 26.025 -12.225 26.195 -4.185 ;
        RECT 26.505 -12.225 26.675 -4.185 ;
        RECT 26.985 -12.225 27.155 -4.185 ;
        RECT 27.465 -12.225 27.635 -4.185 ;
        RECT 27.945 -12.225 28.115 -4.185 ;
        RECT 28.425 -12.225 28.595 -4.185 ;
        RECT 28.905 -12.225 29.075 -4.185 ;
        RECT 29.385 -12.225 29.555 -4.185 ;
        RECT 29.865 -12.225 30.035 -4.185 ;
        RECT 30.345 -12.225 30.515 -4.185 ;
        RECT 30.825 -12.225 30.995 -4.185 ;
        RECT 31.305 -12.225 31.475 -4.185 ;
        RECT 31.785 -12.225 31.955 -4.185 ;
        RECT 32.265 -12.225 32.435 -4.185 ;
        RECT 32.745 -12.225 32.915 -4.185 ;
        RECT 33.225 -12.225 33.395 -4.185 ;
        RECT 33.705 -12.225 33.875 -4.185 ;
        RECT 34.185 -12.225 34.355 -4.185 ;
        RECT 34.665 -12.225 34.835 -4.185 ;
        RECT 35.145 -12.225 35.315 -4.185 ;
        RECT 35.625 -12.225 35.795 -4.185 ;
        RECT 36.105 -12.225 36.275 -4.185 ;
        RECT 36.585 -12.225 36.755 -4.185 ;
        RECT 37.065 -12.225 37.235 -4.185 ;
        RECT 37.545 -12.225 37.715 -4.185 ;
        RECT 38.025 -12.225 38.195 -4.185 ;
        RECT 38.505 -12.225 38.675 -4.185 ;
        RECT 38.985 -12.225 39.155 -4.185 ;
        RECT 39.465 -12.225 39.635 -4.185 ;
        RECT 39.935 -12.225 40.105 -4.185 ;
        RECT 40.415 -12.225 40.585 -4.185 ;
        RECT 40.895 -12.225 41.065 -4.185 ;
        RECT 41.375 -12.225 41.545 -4.185 ;
        RECT 41.855 -12.225 42.025 -4.185 ;
        RECT 42.335 -12.225 42.505 -4.185 ;
        RECT 42.815 -12.225 42.985 -4.185 ;
        RECT 43.295 -12.225 43.465 -4.185 ;
        RECT 43.775 -12.225 43.945 -4.185 ;
        RECT 44.255 -12.225 44.425 -4.185 ;
        RECT 44.735 -12.225 44.905 -4.185 ;
        RECT 45.215 -12.225 45.385 -4.185 ;
        RECT 45.695 -12.225 45.865 -4.185 ;
        RECT 46.175 -12.225 46.345 -4.185 ;
        RECT 46.655 -12.225 46.825 -4.185 ;
        RECT 47.135 -12.225 47.305 -4.185 ;
        RECT 47.615 -12.225 47.785 -4.185 ;
        RECT 48.095 -12.225 48.265 -4.185 ;
        RECT 48.575 -12.225 48.745 -4.185 ;
        RECT 49.055 -12.225 49.225 -4.185 ;
        RECT 49.535 -12.225 49.705 -4.185 ;
        RECT 50.015 -12.225 50.185 -4.185 ;
        RECT 50.495 -12.225 50.665 -4.185 ;
        RECT 50.975 -12.225 51.145 -4.185 ;
        RECT 51.455 -12.225 51.625 -4.185 ;
        RECT 51.935 -12.225 52.105 -4.185 ;
        RECT 52.415 -12.225 52.585 -4.185 ;
        RECT 52.895 -12.225 53.065 -4.185 ;
        RECT 53.375 -12.225 53.545 -4.185 ;
        RECT 53.855 -12.225 54.025 -4.185 ;
        RECT 54.335 -12.225 54.505 -4.185 ;
        RECT 54.815 -12.225 54.985 -4.185 ;
        RECT 55.295 -12.225 55.465 -4.185 ;
        RECT 55.775 -12.225 55.945 -4.185 ;
        RECT 56.255 -12.225 56.425 -4.185 ;
        RECT 56.735 -12.225 56.905 -4.185 ;
        RECT 57.215 -12.225 57.385 -4.185 ;
        RECT 57.695 -12.225 57.865 -4.185 ;
        RECT 58.175 -12.225 58.345 -4.185 ;
        RECT 58.655 -12.225 58.825 -4.185 ;
        RECT 59.135 -12.225 59.305 -4.185 ;
        RECT 59.615 -12.225 59.785 -4.185 ;
        RECT 60.095 -12.225 60.265 -4.185 ;
        RECT 60.575 -12.225 60.745 -4.185 ;
        RECT 61.055 -12.225 61.225 -4.185 ;
        RECT 61.535 -12.225 61.705 -4.185 ;
        RECT 62.015 -12.225 62.185 -4.185 ;
        RECT 62.495 -12.225 62.665 -4.185 ;
        RECT 62.975 -12.225 63.145 -4.185 ;
        RECT 63.455 -12.225 63.625 -4.185 ;
        RECT 63.935 -12.225 64.105 -4.185 ;
        RECT 64.415 -12.225 64.585 -4.185 ;
        RECT 64.895 -12.225 65.065 -4.185 ;
        RECT 65.375 -12.225 65.545 -4.185 ;
        RECT 65.855 -12.225 66.025 -4.185 ;
        RECT 66.335 -12.225 66.505 -4.185 ;
        RECT 66.815 -12.225 66.985 -4.185 ;
        RECT 67.295 -12.225 67.465 -4.185 ;
        RECT 67.775 -12.225 67.945 -4.185 ;
        RECT 68.255 -12.225 68.425 -4.185 ;
        RECT 9.570 -12.230 10.265 -12.225 ;
        RECT 9.235 -12.645 9.565 -12.415 ;
        RECT 10.095 -12.945 10.265 -12.230 ;
        RECT 10.825 -12.625 11.155 -12.455 ;
        RECT 11.785 -12.625 12.115 -12.455 ;
        RECT 12.745 -12.625 13.075 -12.455 ;
        RECT 13.705 -12.625 14.035 -12.455 ;
        RECT 14.665 -12.625 14.995 -12.455 ;
        RECT 15.625 -12.625 15.955 -12.455 ;
        RECT 16.585 -12.625 16.915 -12.455 ;
        RECT 17.545 -12.625 17.875 -12.455 ;
        RECT 18.505 -12.625 18.835 -12.455 ;
        RECT 19.465 -12.625 19.795 -12.455 ;
        RECT 20.425 -12.625 20.755 -12.455 ;
        RECT 21.385 -12.625 21.715 -12.455 ;
        RECT 22.345 -12.625 22.675 -12.455 ;
        RECT 23.305 -12.625 23.635 -12.455 ;
        RECT 24.265 -12.625 24.595 -12.455 ;
        RECT 25.225 -12.625 25.555 -12.455 ;
        RECT 26.185 -12.625 26.515 -12.455 ;
        RECT 27.145 -12.625 27.475 -12.455 ;
        RECT 28.105 -12.615 28.435 -12.445 ;
        RECT 29.065 -12.615 29.395 -12.445 ;
        RECT 30.025 -12.615 30.355 -12.445 ;
        RECT 30.985 -12.615 31.315 -12.445 ;
        RECT 31.945 -12.615 32.275 -12.445 ;
        RECT 32.905 -12.615 33.235 -12.445 ;
        RECT 33.865 -12.615 34.195 -12.445 ;
        RECT 34.825 -12.615 35.155 -12.445 ;
        RECT 35.785 -12.615 36.115 -12.445 ;
        RECT 36.745 -12.615 37.075 -12.445 ;
        RECT 37.705 -12.615 38.035 -12.445 ;
        RECT 38.665 -12.615 38.995 -12.445 ;
        RECT 39.615 -12.615 39.945 -12.445 ;
        RECT 40.575 -12.615 40.905 -12.445 ;
        RECT 41.535 -12.615 41.865 -12.445 ;
        RECT 42.495 -12.615 42.825 -12.445 ;
        RECT 43.455 -12.615 43.785 -12.445 ;
        RECT 44.415 -12.615 44.745 -12.445 ;
        RECT 45.375 -12.615 45.705 -12.445 ;
        RECT 46.335 -12.615 46.665 -12.445 ;
        RECT 47.295 -12.615 47.625 -12.445 ;
        RECT 48.255 -12.615 48.585 -12.445 ;
        RECT 49.215 -12.615 49.545 -12.445 ;
        RECT 50.175 -12.615 50.505 -12.445 ;
        RECT 51.135 -12.615 51.465 -12.445 ;
        RECT 52.095 -12.615 52.425 -12.445 ;
        RECT 53.055 -12.615 53.385 -12.445 ;
        RECT 54.015 -12.615 54.345 -12.445 ;
        RECT 54.975 -12.615 55.305 -12.445 ;
        RECT 55.935 -12.615 56.265 -12.445 ;
        RECT 56.895 -12.615 57.225 -12.445 ;
        RECT 57.855 -12.615 58.185 -12.445 ;
        RECT 58.815 -12.615 59.145 -12.445 ;
        RECT 59.775 -12.615 60.105 -12.445 ;
        RECT 60.735 -12.615 61.065 -12.445 ;
        RECT 61.695 -12.615 62.025 -12.445 ;
        RECT 62.655 -12.615 62.985 -12.445 ;
        RECT 63.615 -12.615 63.945 -12.445 ;
        RECT 64.575 -12.615 64.905 -12.445 ;
        RECT 65.535 -12.615 65.865 -12.445 ;
        RECT 66.495 -12.615 66.825 -12.445 ;
        RECT 67.455 -12.615 67.785 -12.445 ;
        RECT 68.825 -12.945 68.995 -3.470 ;
        RECT 8.525 -13.115 68.995 -12.945 ;
      LAYER met1 ;
        RECT 5.520 106.300 167.900 106.470 ;
        RECT 167.990 106.300 168.570 106.470 ;
        RECT 5.520 106.130 168.570 106.300 ;
        RECT 5.520 0.000 167.900 106.130 ;
        RECT 167.990 105.960 168.570 106.130 ;
        RECT 8.620 -3.500 68.900 -3.260 ;
        RECT 8.630 -3.580 68.890 -3.500 ;
        RECT 9.810 -3.600 68.890 -3.580 ;
        RECT 9.165 -3.770 9.625 -3.735 ;
        RECT 7.130 -3.810 9.625 -3.770 ;
        RECT 7.065 -3.890 9.625 -3.810 ;
        RECT 7.065 -4.040 9.630 -3.890 ;
        RECT 10.100 -4.000 68.250 -3.760 ;
        RECT 6.370 -9.110 6.750 -9.050 ;
        RECT 6.350 -11.250 6.770 -9.110 ;
        RECT 6.370 -11.310 6.750 -11.250 ;
        RECT 6.925 -12.200 7.155 -4.200 ;
        RECT 7.395 -4.205 9.170 -4.200 ;
        RECT 7.395 -12.200 9.295 -4.205 ;
        RECT 9.065 -12.205 9.295 -12.200 ;
        RECT 9.505 -12.205 9.735 -4.205 ;
        RECT 10.100 -7.550 10.340 -4.000 ;
        RECT 9.880 -8.790 10.390 -7.550 ;
        RECT 7.055 -12.415 9.530 -12.360 ;
        RECT 10.100 -12.410 10.340 -8.790 ;
        RECT 10.635 -9.210 10.865 -4.205 ;
        RECT 11.030 -7.200 11.420 -4.200 ;
        RECT 10.550 -12.210 10.940 -9.210 ;
        RECT 11.115 -12.205 11.345 -7.200 ;
        RECT 11.595 -9.210 11.825 -4.205 ;
        RECT 11.990 -7.200 12.380 -4.200 ;
        RECT 11.510 -12.210 11.900 -9.210 ;
        RECT 12.075 -12.205 12.305 -7.200 ;
        RECT 12.555 -9.210 12.785 -4.205 ;
        RECT 12.950 -7.200 13.340 -4.200 ;
        RECT 12.470 -12.210 12.860 -9.210 ;
        RECT 13.035 -12.205 13.265 -7.200 ;
        RECT 13.515 -9.210 13.745 -4.205 ;
        RECT 13.910 -7.200 14.300 -4.200 ;
        RECT 13.430 -12.210 13.820 -9.210 ;
        RECT 13.995 -12.205 14.225 -7.200 ;
        RECT 14.475 -9.210 14.705 -4.205 ;
        RECT 14.870 -7.200 15.260 -4.200 ;
        RECT 14.390 -12.210 14.780 -9.210 ;
        RECT 14.955 -12.205 15.185 -7.200 ;
        RECT 15.435 -9.210 15.665 -4.205 ;
        RECT 15.830 -7.200 16.220 -4.200 ;
        RECT 15.350 -12.210 15.740 -9.210 ;
        RECT 15.915 -12.205 16.145 -7.200 ;
        RECT 16.395 -9.210 16.625 -4.205 ;
        RECT 16.790 -7.200 17.180 -4.200 ;
        RECT 16.310 -12.210 16.700 -9.210 ;
        RECT 16.875 -12.205 17.105 -7.200 ;
        RECT 17.355 -9.210 17.585 -4.205 ;
        RECT 17.750 -7.200 18.140 -4.200 ;
        RECT 17.270 -12.210 17.660 -9.210 ;
        RECT 17.835 -12.205 18.065 -7.200 ;
        RECT 18.315 -9.210 18.545 -4.205 ;
        RECT 18.710 -7.200 19.100 -4.200 ;
        RECT 18.230 -12.210 18.620 -9.210 ;
        RECT 18.795 -12.205 19.025 -7.200 ;
        RECT 19.275 -9.210 19.505 -4.205 ;
        RECT 19.755 -4.210 19.985 -4.205 ;
        RECT 19.670 -7.210 20.060 -4.210 ;
        RECT 19.190 -12.210 19.580 -9.210 ;
        RECT 19.755 -12.205 19.985 -7.210 ;
        RECT 20.235 -9.210 20.465 -4.205 ;
        RECT 20.715 -4.210 20.945 -4.205 ;
        RECT 20.630 -7.210 21.020 -4.210 ;
        RECT 20.150 -12.210 20.540 -9.210 ;
        RECT 20.715 -12.205 20.945 -7.210 ;
        RECT 21.195 -9.210 21.425 -4.205 ;
        RECT 21.675 -4.210 21.905 -4.205 ;
        RECT 21.590 -7.210 21.980 -4.210 ;
        RECT 21.110 -12.210 21.500 -9.210 ;
        RECT 21.675 -12.205 21.905 -7.210 ;
        RECT 22.155 -9.210 22.385 -4.205 ;
        RECT 22.635 -4.210 22.865 -4.205 ;
        RECT 22.550 -7.210 22.940 -4.210 ;
        RECT 22.070 -12.210 22.460 -9.210 ;
        RECT 22.635 -12.205 22.865 -7.210 ;
        RECT 23.115 -9.210 23.345 -4.205 ;
        RECT 23.595 -4.210 23.825 -4.205 ;
        RECT 23.510 -7.210 23.900 -4.210 ;
        RECT 23.030 -12.210 23.420 -9.210 ;
        RECT 23.595 -12.205 23.825 -7.210 ;
        RECT 24.075 -9.210 24.305 -4.205 ;
        RECT 24.555 -4.210 24.785 -4.205 ;
        RECT 24.470 -7.210 24.860 -4.210 ;
        RECT 23.990 -12.210 24.380 -9.210 ;
        RECT 24.555 -12.205 24.785 -7.210 ;
        RECT 25.035 -9.210 25.265 -4.205 ;
        RECT 25.515 -4.210 25.745 -4.205 ;
        RECT 25.430 -7.210 25.820 -4.210 ;
        RECT 24.950 -12.210 25.340 -9.210 ;
        RECT 25.515 -12.205 25.745 -7.210 ;
        RECT 25.995 -9.210 26.225 -4.205 ;
        RECT 26.475 -4.210 26.705 -4.205 ;
        RECT 26.390 -7.210 26.780 -4.210 ;
        RECT 25.910 -12.210 26.300 -9.210 ;
        RECT 26.475 -12.205 26.705 -7.210 ;
        RECT 26.955 -9.210 27.185 -4.205 ;
        RECT 27.435 -4.210 27.665 -4.205 ;
        RECT 27.350 -7.210 27.740 -4.210 ;
        RECT 26.870 -12.210 27.260 -9.210 ;
        RECT 27.435 -12.205 27.665 -7.210 ;
        RECT 27.915 -9.210 28.145 -4.205 ;
        RECT 28.395 -4.210 28.625 -4.205 ;
        RECT 28.310 -7.210 28.700 -4.210 ;
        RECT 27.830 -12.210 28.220 -9.210 ;
        RECT 28.395 -12.205 28.625 -7.210 ;
        RECT 28.875 -9.210 29.105 -4.205 ;
        RECT 29.355 -4.210 29.585 -4.205 ;
        RECT 29.270 -7.210 29.660 -4.210 ;
        RECT 28.790 -12.210 29.180 -9.210 ;
        RECT 29.355 -12.205 29.585 -7.210 ;
        RECT 29.835 -9.210 30.065 -4.205 ;
        RECT 30.315 -4.210 30.545 -4.205 ;
        RECT 30.230 -7.210 30.620 -4.210 ;
        RECT 29.750 -12.210 30.140 -9.210 ;
        RECT 30.315 -12.205 30.545 -7.210 ;
        RECT 30.795 -9.210 31.025 -4.205 ;
        RECT 31.275 -4.210 31.505 -4.205 ;
        RECT 31.190 -7.210 31.580 -4.210 ;
        RECT 30.710 -12.210 31.100 -9.210 ;
        RECT 31.275 -12.205 31.505 -7.210 ;
        RECT 31.755 -9.210 31.985 -4.205 ;
        RECT 32.235 -4.210 32.465 -4.205 ;
        RECT 32.150 -7.210 32.540 -4.210 ;
        RECT 31.670 -12.210 32.060 -9.210 ;
        RECT 32.235 -12.205 32.465 -7.210 ;
        RECT 32.715 -9.210 32.945 -4.205 ;
        RECT 33.195 -4.210 33.425 -4.205 ;
        RECT 33.110 -7.210 33.500 -4.210 ;
        RECT 32.630 -12.210 33.020 -9.210 ;
        RECT 33.195 -12.205 33.425 -7.210 ;
        RECT 33.675 -9.210 33.905 -4.205 ;
        RECT 34.155 -4.210 34.385 -4.205 ;
        RECT 34.070 -7.210 34.460 -4.210 ;
        RECT 33.590 -12.210 33.980 -9.210 ;
        RECT 34.155 -12.205 34.385 -7.210 ;
        RECT 34.635 -9.210 34.865 -4.205 ;
        RECT 35.115 -4.210 35.345 -4.205 ;
        RECT 35.030 -7.210 35.420 -4.210 ;
        RECT 34.550 -12.210 34.940 -9.210 ;
        RECT 35.115 -12.205 35.345 -7.210 ;
        RECT 35.595 -9.210 35.825 -4.205 ;
        RECT 36.075 -4.210 36.305 -4.205 ;
        RECT 35.990 -7.210 36.380 -4.210 ;
        RECT 35.510 -12.210 35.900 -9.210 ;
        RECT 36.075 -12.205 36.305 -7.210 ;
        RECT 36.555 -9.210 36.785 -4.205 ;
        RECT 37.035 -4.210 37.265 -4.205 ;
        RECT 36.950 -7.210 37.340 -4.210 ;
        RECT 36.470 -12.210 36.860 -9.210 ;
        RECT 37.035 -12.205 37.265 -7.210 ;
        RECT 37.515 -9.210 37.745 -4.205 ;
        RECT 37.995 -4.210 38.225 -4.205 ;
        RECT 37.910 -7.210 38.300 -4.210 ;
        RECT 37.430 -12.210 37.820 -9.210 ;
        RECT 37.995 -12.205 38.225 -7.210 ;
        RECT 38.475 -9.210 38.705 -4.205 ;
        RECT 38.955 -4.210 39.185 -4.205 ;
        RECT 38.870 -7.210 39.260 -4.210 ;
        RECT 38.390 -12.210 38.780 -9.210 ;
        RECT 38.955 -12.205 39.185 -7.210 ;
        RECT 39.435 -9.210 39.665 -4.205 ;
        RECT 39.905 -4.210 40.135 -4.205 ;
        RECT 39.830 -7.210 40.220 -4.210 ;
        RECT 39.350 -12.210 39.740 -9.210 ;
        RECT 39.905 -12.205 40.135 -7.210 ;
        RECT 40.385 -9.210 40.615 -4.205 ;
        RECT 40.865 -4.210 41.095 -4.205 ;
        RECT 40.790 -7.210 41.180 -4.210 ;
        RECT 40.310 -12.210 40.700 -9.210 ;
        RECT 40.865 -12.205 41.095 -7.210 ;
        RECT 41.345 -9.210 41.575 -4.205 ;
        RECT 41.825 -4.210 42.055 -4.205 ;
        RECT 41.750 -7.210 42.140 -4.210 ;
        RECT 41.270 -12.210 41.660 -9.210 ;
        RECT 41.825 -12.205 42.055 -7.210 ;
        RECT 42.305 -9.210 42.535 -4.205 ;
        RECT 42.785 -4.210 43.015 -4.205 ;
        RECT 42.710 -7.210 43.100 -4.210 ;
        RECT 42.230 -12.210 42.620 -9.210 ;
        RECT 42.785 -12.205 43.015 -7.210 ;
        RECT 43.265 -9.210 43.495 -4.205 ;
        RECT 43.745 -4.210 43.975 -4.205 ;
        RECT 43.670 -7.210 44.060 -4.210 ;
        RECT 43.190 -12.210 43.580 -9.210 ;
        RECT 43.745 -12.205 43.975 -7.210 ;
        RECT 44.225 -9.210 44.455 -4.205 ;
        RECT 44.705 -4.210 44.935 -4.205 ;
        RECT 44.630 -7.210 45.020 -4.210 ;
        RECT 44.150 -12.210 44.540 -9.210 ;
        RECT 44.705 -12.205 44.935 -7.210 ;
        RECT 45.185 -9.210 45.415 -4.205 ;
        RECT 45.665 -4.210 45.895 -4.205 ;
        RECT 45.590 -7.210 45.980 -4.210 ;
        RECT 45.110 -12.210 45.500 -9.210 ;
        RECT 45.665 -12.205 45.895 -7.210 ;
        RECT 46.145 -9.210 46.375 -4.205 ;
        RECT 46.625 -4.210 46.855 -4.205 ;
        RECT 46.550 -7.210 46.940 -4.210 ;
        RECT 46.070 -12.210 46.460 -9.210 ;
        RECT 46.625 -12.205 46.855 -7.210 ;
        RECT 47.105 -9.210 47.335 -4.205 ;
        RECT 47.585 -4.210 47.815 -4.205 ;
        RECT 47.510 -7.210 47.900 -4.210 ;
        RECT 47.030 -12.210 47.420 -9.210 ;
        RECT 47.585 -12.205 47.815 -7.210 ;
        RECT 48.065 -9.210 48.295 -4.205 ;
        RECT 48.545 -4.210 48.775 -4.205 ;
        RECT 48.470 -7.210 48.860 -4.210 ;
        RECT 47.990 -12.210 48.380 -9.210 ;
        RECT 48.545 -12.205 48.775 -7.210 ;
        RECT 49.025 -9.210 49.255 -4.205 ;
        RECT 49.505 -4.210 49.735 -4.205 ;
        RECT 49.430 -7.210 49.820 -4.210 ;
        RECT 48.950 -12.210 49.340 -9.210 ;
        RECT 49.505 -12.205 49.735 -7.210 ;
        RECT 49.985 -9.210 50.215 -4.205 ;
        RECT 50.465 -4.210 50.695 -4.205 ;
        RECT 50.390 -7.210 50.780 -4.210 ;
        RECT 49.910 -12.210 50.300 -9.210 ;
        RECT 50.465 -12.205 50.695 -7.210 ;
        RECT 50.945 -9.210 51.175 -4.205 ;
        RECT 51.425 -4.210 51.655 -4.205 ;
        RECT 51.350 -7.210 51.740 -4.210 ;
        RECT 50.870 -12.210 51.260 -9.210 ;
        RECT 51.425 -12.205 51.655 -7.210 ;
        RECT 51.905 -9.210 52.135 -4.205 ;
        RECT 52.385 -4.210 52.615 -4.205 ;
        RECT 52.310 -7.210 52.700 -4.210 ;
        RECT 51.830 -12.210 52.220 -9.210 ;
        RECT 52.385 -12.205 52.615 -7.210 ;
        RECT 52.865 -9.210 53.095 -4.205 ;
        RECT 53.345 -4.210 53.575 -4.205 ;
        RECT 53.270 -7.210 53.660 -4.210 ;
        RECT 52.790 -12.210 53.180 -9.210 ;
        RECT 53.345 -12.205 53.575 -7.210 ;
        RECT 53.825 -9.210 54.055 -4.205 ;
        RECT 54.305 -4.210 54.535 -4.205 ;
        RECT 54.230 -7.210 54.620 -4.210 ;
        RECT 53.750 -12.210 54.140 -9.210 ;
        RECT 54.305 -12.205 54.535 -7.210 ;
        RECT 54.785 -9.210 55.015 -4.205 ;
        RECT 55.265 -4.210 55.495 -4.205 ;
        RECT 55.190 -7.210 55.580 -4.210 ;
        RECT 54.710 -12.210 55.100 -9.210 ;
        RECT 55.265 -12.205 55.495 -7.210 ;
        RECT 55.745 -9.210 55.975 -4.205 ;
        RECT 56.225 -4.210 56.455 -4.205 ;
        RECT 56.150 -7.210 56.540 -4.210 ;
        RECT 55.670 -12.210 56.060 -9.210 ;
        RECT 56.225 -12.205 56.455 -7.210 ;
        RECT 56.705 -9.210 56.935 -4.205 ;
        RECT 57.185 -4.210 57.415 -4.205 ;
        RECT 57.110 -7.210 57.500 -4.210 ;
        RECT 56.630 -12.210 57.020 -9.210 ;
        RECT 57.185 -12.205 57.415 -7.210 ;
        RECT 57.665 -9.210 57.895 -4.205 ;
        RECT 58.145 -4.210 58.375 -4.205 ;
        RECT 58.070 -7.210 58.460 -4.210 ;
        RECT 57.590 -12.210 57.980 -9.210 ;
        RECT 58.145 -12.205 58.375 -7.210 ;
        RECT 58.625 -9.210 58.855 -4.205 ;
        RECT 59.105 -4.210 59.335 -4.205 ;
        RECT 59.030 -7.210 59.420 -4.210 ;
        RECT 58.550 -12.210 58.940 -9.210 ;
        RECT 59.105 -12.205 59.335 -7.210 ;
        RECT 59.585 -9.210 59.815 -4.205 ;
        RECT 60.065 -4.210 60.295 -4.205 ;
        RECT 59.990 -7.210 60.380 -4.210 ;
        RECT 59.510 -12.210 59.900 -9.210 ;
        RECT 60.065 -12.205 60.295 -7.210 ;
        RECT 60.545 -9.210 60.775 -4.205 ;
        RECT 61.025 -4.210 61.255 -4.205 ;
        RECT 60.950 -7.210 61.340 -4.210 ;
        RECT 60.470 -12.210 60.860 -9.210 ;
        RECT 61.025 -12.205 61.255 -7.210 ;
        RECT 61.505 -9.210 61.735 -4.205 ;
        RECT 61.985 -4.210 62.215 -4.205 ;
        RECT 61.910 -7.210 62.300 -4.210 ;
        RECT 61.430 -12.210 61.820 -9.210 ;
        RECT 61.985 -12.205 62.215 -7.210 ;
        RECT 62.465 -9.210 62.695 -4.205 ;
        RECT 62.945 -4.210 63.175 -4.205 ;
        RECT 62.870 -7.210 63.260 -4.210 ;
        RECT 62.390 -12.210 62.780 -9.210 ;
        RECT 62.945 -12.205 63.175 -7.210 ;
        RECT 63.425 -9.210 63.655 -4.205 ;
        RECT 63.905 -4.210 64.135 -4.205 ;
        RECT 63.830 -7.210 64.220 -4.210 ;
        RECT 63.350 -12.210 63.740 -9.210 ;
        RECT 63.905 -12.205 64.135 -7.210 ;
        RECT 64.385 -9.210 64.615 -4.205 ;
        RECT 64.865 -4.210 65.095 -4.205 ;
        RECT 64.790 -7.210 65.180 -4.210 ;
        RECT 64.310 -12.210 64.700 -9.210 ;
        RECT 64.865 -12.205 65.095 -7.210 ;
        RECT 65.345 -9.210 65.575 -4.205 ;
        RECT 65.825 -4.210 66.055 -4.205 ;
        RECT 65.750 -7.210 66.140 -4.210 ;
        RECT 65.270 -12.210 65.660 -9.210 ;
        RECT 65.825 -12.205 66.055 -7.210 ;
        RECT 66.305 -9.210 66.535 -4.205 ;
        RECT 66.785 -4.210 67.015 -4.205 ;
        RECT 66.710 -7.210 67.100 -4.210 ;
        RECT 66.230 -12.210 66.620 -9.210 ;
        RECT 66.785 -12.205 67.015 -7.210 ;
        RECT 67.265 -9.210 67.495 -4.205 ;
        RECT 67.745 -4.210 67.975 -4.205 ;
        RECT 67.670 -7.210 68.060 -4.210 ;
        RECT 67.190 -12.210 67.580 -9.210 ;
        RECT 67.745 -12.205 67.975 -7.210 ;
        RECT 68.225 -9.210 68.455 -4.205 ;
        RECT 68.150 -12.210 68.540 -9.210 ;
        RECT 7.055 -12.590 9.615 -12.415 ;
        RECT 7.070 -12.650 9.615 -12.590 ;
        RECT 10.100 -12.650 67.770 -12.410 ;
        RECT 9.155 -12.665 9.615 -12.650 ;
        RECT 10.845 -12.655 11.135 -12.650 ;
        RECT 11.805 -12.655 12.095 -12.650 ;
        RECT 12.765 -12.655 13.055 -12.650 ;
        RECT 13.725 -12.655 14.015 -12.650 ;
        RECT 14.685 -12.655 14.975 -12.650 ;
        RECT 15.645 -12.655 15.935 -12.650 ;
        RECT 16.605 -12.655 16.895 -12.650 ;
        RECT 17.565 -12.655 17.855 -12.650 ;
        RECT 18.525 -12.655 18.815 -12.650 ;
        RECT 19.485 -12.655 19.775 -12.650 ;
        RECT 20.445 -12.655 20.735 -12.650 ;
        RECT 21.405 -12.655 21.695 -12.650 ;
        RECT 22.365 -12.655 22.655 -12.650 ;
        RECT 23.325 -12.655 23.615 -12.650 ;
        RECT 24.285 -12.655 24.575 -12.650 ;
        RECT 25.245 -12.655 25.535 -12.650 ;
        RECT 26.205 -12.655 26.495 -12.650 ;
        RECT 27.165 -12.655 27.455 -12.650 ;
      LAYER met2 ;
        RECT 6.270 0.000 167.900 107.285 ;
        RECT 167.990 105.960 168.570 106.470 ;
        RECT 8.680 -3.650 68.840 -3.240 ;
        RECT 11.080 -7.300 68.020 -4.110 ;
        RECT 8.460 -8.840 10.340 -7.490 ;
        RECT 6.400 -11.300 6.720 -9.060 ;
        RECT 6.270 -12.800 7.880 -12.210 ;
        RECT 10.600 -12.310 68.490 -9.110 ;
      LAYER met3 ;
        RECT 1.300 0.000 167.900 107.265 ;
        RECT 167.990 105.960 168.570 106.470 ;
        RECT 6.210 -7.250 69.180 -3.110 ;
        RECT 11.030 -7.275 69.180 -7.250 ;
        RECT 68.020 -7.280 69.180 -7.275 ;
        RECT 6.350 -9.100 6.770 -9.085 ;
        RECT 1.300 -9.110 6.830 -9.100 ;
        RECT 1.300 -11.200 7.910 -9.110 ;
        RECT 1.300 -16.440 3.400 -11.200 ;
        RECT 6.220 -11.260 7.910 -11.200 ;
        RECT 6.350 -11.275 6.770 -11.260 ;
        RECT 6.220 -13.320 7.910 -12.230 ;
        RECT 8.320 -13.320 69.190 -9.110 ;
        RECT 91.260 -16.440 94.780 -15.890 ;
        RECT 1.300 -18.540 94.780 -16.440 ;
        RECT 91.260 -19.050 94.780 -18.540 ;
      LAYER met4 ;
        RECT 1.210 103.530 7.270 108.100 ;
        RECT 1.210 100.330 1.250 103.130 ;
        RECT 3.175 100.060 7.270 103.530 ;
        RECT 8.370 102.100 10.950 108.100 ;
        RECT 12.050 102.100 14.630 108.100 ;
        RECT 15.730 102.100 18.310 108.100 ;
        RECT 19.410 102.100 21.990 108.100 ;
        RECT 23.090 104.140 25.670 108.100 ;
        RECT 26.770 104.140 29.350 108.100 ;
        RECT 23.090 102.100 29.350 104.140 ;
        RECT 30.450 102.100 33.030 108.100 ;
        RECT 8.370 100.060 33.030 102.100 ;
        RECT 34.130 100.060 36.710 108.100 ;
        RECT 37.810 100.060 40.390 108.100 ;
        RECT 41.490 106.860 44.070 108.100 ;
        RECT 45.170 106.860 47.750 108.100 ;
        RECT 48.850 106.860 51.430 108.100 ;
        RECT 41.490 104.000 51.430 106.860 ;
        RECT 41.490 100.060 43.530 104.000 ;
        RECT 3.175 4.800 43.530 100.060 ;
        RECT 45.930 100.060 51.430 104.000 ;
        RECT 52.530 106.860 55.110 108.100 ;
        RECT 56.210 106.860 58.790 108.100 ;
        RECT 59.890 106.860 62.470 108.100 ;
        RECT 52.530 101.420 62.470 106.860 ;
        RECT 63.570 106.860 66.150 108.100 ;
        RECT 67.250 106.860 69.830 108.100 ;
        RECT 63.570 106.180 69.830 106.860 ;
        RECT 70.930 106.860 73.510 108.100 ;
        RECT 74.610 106.860 77.190 108.100 ;
        RECT 78.290 106.860 80.870 108.100 ;
        RECT 81.970 106.860 84.550 108.100 ;
        RECT 70.930 106.180 84.550 106.860 ;
        RECT 85.650 106.860 88.230 108.100 ;
        RECT 89.330 106.860 91.910 108.100 ;
        RECT 93.010 107.400 95.590 108.100 ;
        RECT 96.690 107.400 99.270 108.100 ;
        RECT 93.010 106.860 99.270 107.400 ;
        RECT 100.370 106.860 102.950 108.100 ;
        RECT 85.650 106.180 102.950 106.860 ;
        RECT 63.570 104.140 102.950 106.180 ;
        RECT 104.050 106.860 106.630 108.100 ;
        RECT 107.730 106.860 110.310 108.100 ;
        RECT 111.410 106.860 113.990 108.100 ;
        RECT 104.050 104.140 113.990 106.860 ;
        RECT 63.570 104.000 113.990 104.140 ;
        RECT 63.570 101.420 82.740 104.000 ;
        RECT 52.530 100.060 82.740 101.420 ;
        RECT 45.930 4.800 82.740 100.060 ;
        RECT 85.140 102.100 113.990 104.000 ;
        RECT 115.090 106.860 117.670 108.100 ;
        RECT 118.770 106.860 121.350 108.100 ;
        RECT 122.450 107.400 125.030 108.100 ;
        RECT 126.130 107.400 128.710 108.100 ;
        RECT 122.450 106.860 128.710 107.400 ;
        RECT 129.810 106.860 132.390 108.100 ;
        RECT 115.090 104.820 132.390 106.860 ;
        RECT 133.490 106.860 136.070 108.100 ;
        RECT 137.170 106.860 139.750 108.100 ;
        RECT 133.490 104.820 139.750 106.860 ;
        RECT 140.850 106.860 143.430 108.100 ;
        RECT 144.530 106.860 147.110 108.100 ;
        RECT 140.850 104.820 147.110 106.860 ;
        RECT 148.210 106.860 150.790 108.100 ;
        RECT 151.890 107.400 154.470 108.100 ;
        RECT 155.570 107.400 158.150 108.100 ;
        RECT 159.250 107.400 161.830 108.100 ;
        RECT 162.930 107.400 167.900 108.100 ;
        RECT 151.890 106.860 167.900 107.400 ;
        RECT 148.210 104.820 167.900 106.860 ;
        RECT 167.990 106.150 168.570 106.470 ;
        RECT 167.990 105.700 168.580 106.150 ;
        RECT 168.020 105.080 168.580 105.700 ;
        RECT 115.090 104.000 167.900 104.820 ;
        RECT 115.090 102.100 121.950 104.000 ;
        RECT 85.140 4.800 121.950 102.100 ;
        RECT 124.350 4.800 161.160 104.000 ;
        RECT 161.560 4.800 163.160 5.200 ;
        RECT 163.560 4.800 167.900 104.000 ;
        RECT 3.175 0.000 167.900 4.800 ;
        RECT 2.775 -2.010 12.180 -0.485 ;
        RECT 10.660 -3.025 12.170 -2.010 ;
        RECT 10.660 -4.535 68.985 -3.025 ;
        RECT 79.410 -11.600 81.010 0.000 ;
        RECT 161.560 -0.700 163.160 0.000 ;
        RECT 5.290 -15.160 7.840 -12.230 ;
        RECT 10.600 -13.200 81.010 -11.600 ;
        RECT 92.650 -2.300 163.160 -0.700 ;
        RECT 5.790 -21.390 6.370 -15.160 ;
        RECT 92.650 -15.890 94.250 -2.300 ;
        RECT 101.340 -8.525 101.920 -8.510 ;
        RECT 168.025 -8.525 168.575 105.080 ;
        RECT 101.340 -9.075 168.575 -8.525 ;
        RECT 91.260 -19.050 94.780 -15.890 ;
        RECT 101.340 -21.390 101.920 -9.075 ;
        RECT 5.790 -21.970 101.920 -21.390 ;
  END
END tt_um_power_test
END LIBRARY

