VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_test
  CLASS BLOCK ;
  FOREIGN tt_um_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 106.950 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 107.260 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 107.260 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 107.800 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 107.800 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 107.800 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 107.800 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 107.800 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 107.800 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 107.800 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 107.260 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 102.500 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 107.260 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 107.260 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 107.260 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 107.260 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 107.260 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 107.260 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 100.460 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 100.460 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 104.540 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 100.460 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 97.740 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 100.460 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 100.460 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 97.740 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 102.500 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 100.460 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 106.580 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 107.260 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 97.740 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 107.260 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 107.260 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 107.260 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 103.180 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 107.260 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 104.540 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 103.180 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 107.260 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 103.180 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 107.260 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 107.260 66.850 108.800 ;
    END
  END uo_out[7]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.930 5.200 45.530 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.140 5.200 84.740 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.350 5.200 123.950 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 161.560 5.200 163.160 103.600 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -5.420 -25.800 -0.420 77.240 ;
    END
  END vccd1
  OBS
      LAYER nwell ;
        RECT 17.145 -24.585 34.615 -12.395 ;
      LAYER li1 ;
        RECT 5.520 0.000 162.380 103.445 ;
        RECT 17.325 -12.745 34.435 -12.575 ;
        RECT 17.325 -24.235 17.495 -12.745 ;
        RECT 18.125 -13.255 18.625 -13.085 ;
        RECT 18.915 -13.255 19.415 -13.085 ;
        RECT 19.705 -13.255 20.205 -13.085 ;
        RECT 20.495 -13.255 20.995 -13.085 ;
        RECT 21.285 -13.255 21.785 -13.085 ;
        RECT 22.075 -13.255 22.575 -13.085 ;
        RECT 22.865 -13.255 23.365 -13.085 ;
        RECT 23.655 -13.255 24.155 -13.085 ;
        RECT 24.445 -13.255 24.945 -13.085 ;
        RECT 25.235 -13.255 25.735 -13.085 ;
        RECT 26.025 -13.255 26.525 -13.085 ;
        RECT 26.815 -13.255 27.315 -13.085 ;
        RECT 27.605 -13.255 28.105 -13.085 ;
        RECT 28.395 -13.255 28.895 -13.085 ;
        RECT 29.185 -13.255 29.685 -13.085 ;
        RECT 29.975 -13.255 30.475 -13.085 ;
        RECT 30.765 -13.255 31.265 -13.085 ;
        RECT 31.555 -13.255 32.055 -13.085 ;
        RECT 32.345 -13.255 32.845 -13.085 ;
        RECT 33.135 -13.255 33.635 -13.085 ;
        RECT 17.895 -23.510 18.065 -13.470 ;
        RECT 18.685 -23.510 18.855 -13.470 ;
        RECT 19.475 -23.510 19.645 -13.470 ;
        RECT 20.265 -23.510 20.435 -13.470 ;
        RECT 21.055 -23.510 21.225 -13.470 ;
        RECT 21.845 -23.510 22.015 -13.470 ;
        RECT 22.635 -23.510 22.805 -13.470 ;
        RECT 23.425 -23.510 23.595 -13.470 ;
        RECT 24.215 -23.510 24.385 -13.470 ;
        RECT 25.005 -23.510 25.175 -13.470 ;
        RECT 25.795 -23.510 25.965 -13.470 ;
        RECT 26.585 -23.510 26.755 -13.470 ;
        RECT 27.375 -23.510 27.545 -13.470 ;
        RECT 28.165 -23.510 28.335 -13.470 ;
        RECT 28.955 -23.510 29.125 -13.470 ;
        RECT 29.745 -23.510 29.915 -13.470 ;
        RECT 30.535 -23.510 30.705 -13.470 ;
        RECT 31.325 -23.510 31.495 -13.470 ;
        RECT 32.115 -23.510 32.285 -13.470 ;
        RECT 32.905 -23.510 33.075 -13.470 ;
        RECT 33.695 -23.510 33.865 -13.470 ;
        RECT 18.125 -23.895 18.625 -23.725 ;
        RECT 18.915 -23.895 19.415 -23.725 ;
        RECT 19.705 -23.895 20.205 -23.725 ;
        RECT 20.495 -23.895 20.995 -23.725 ;
        RECT 21.285 -23.895 21.785 -23.725 ;
        RECT 22.075 -23.895 22.575 -23.725 ;
        RECT 22.865 -23.895 23.365 -23.725 ;
        RECT 23.655 -23.895 24.155 -23.725 ;
        RECT 24.445 -23.895 24.945 -23.725 ;
        RECT 25.235 -23.895 25.735 -23.725 ;
        RECT 26.025 -23.895 26.525 -23.725 ;
        RECT 26.815 -23.895 27.315 -23.725 ;
        RECT 27.605 -23.895 28.105 -23.725 ;
        RECT 28.395 -23.895 28.895 -23.725 ;
        RECT 29.185 -23.895 29.685 -23.725 ;
        RECT 29.975 -23.895 30.475 -23.725 ;
        RECT 30.765 -23.895 31.265 -23.725 ;
        RECT 31.555 -23.895 32.055 -23.725 ;
        RECT 32.345 -23.895 32.845 -23.725 ;
        RECT 33.135 -23.895 33.635 -23.725 ;
        RECT 34.265 -24.235 34.435 -12.745 ;
        RECT 17.325 -24.405 34.435 -24.235 ;
      LAYER met1 ;
        RECT 5.520 0.000 163.160 107.060 ;
        RECT 17.820 -12.480 33.950 -12.460 ;
        RECT 35.590 -12.480 37.530 -12.320 ;
        RECT 17.820 -12.490 37.530 -12.480 ;
        RECT 17.680 -12.620 37.530 -12.490 ;
        RECT 14.170 -13.020 15.400 -12.700 ;
        RECT 17.680 -12.780 35.890 -12.620 ;
        RECT 17.680 -12.850 34.130 -12.780 ;
        RECT 14.170 -13.320 33.960 -13.020 ;
        RECT 14.170 -23.660 15.400 -13.320 ;
        RECT 17.865 -13.660 18.095 -13.575 ;
        RECT 19.445 -13.660 19.675 -13.575 ;
        RECT 21.025 -13.660 21.255 -13.575 ;
        RECT 22.605 -13.660 22.835 -13.575 ;
        RECT 24.185 -13.660 24.415 -13.575 ;
        RECT 25.765 -13.660 25.995 -13.575 ;
        RECT 27.345 -13.660 27.575 -13.575 ;
        RECT 28.925 -13.660 29.155 -13.575 ;
        RECT 30.505 -13.660 30.735 -13.575 ;
        RECT 32.085 -13.660 32.315 -13.575 ;
        RECT 33.665 -13.660 33.895 -13.575 ;
        RECT 16.320 -17.970 35.220 -13.660 ;
        RECT 17.865 -18.635 18.095 -17.970 ;
        RECT 18.655 -18.990 18.885 -18.345 ;
        RECT 19.445 -18.635 19.675 -17.970 ;
        RECT 20.235 -18.990 20.465 -18.345 ;
        RECT 21.025 -18.635 21.255 -17.970 ;
        RECT 21.815 -18.990 22.045 -18.345 ;
        RECT 22.605 -18.635 22.835 -17.970 ;
        RECT 23.395 -18.990 23.625 -18.345 ;
        RECT 24.185 -18.635 24.415 -17.970 ;
        RECT 24.975 -18.990 25.205 -18.345 ;
        RECT 25.765 -18.635 25.995 -17.970 ;
        RECT 26.555 -18.990 26.785 -18.345 ;
        RECT 27.345 -18.635 27.575 -17.970 ;
        RECT 28.135 -18.990 28.365 -18.345 ;
        RECT 28.925 -18.635 29.155 -17.970 ;
        RECT 29.715 -18.990 29.945 -18.345 ;
        RECT 30.505 -18.635 30.735 -17.970 ;
        RECT 31.295 -18.990 31.525 -18.345 ;
        RECT 32.085 -18.635 32.315 -17.970 ;
        RECT 32.875 -18.990 33.105 -18.345 ;
        RECT 33.665 -18.635 33.895 -17.970 ;
        RECT 16.340 -23.300 35.240 -18.990 ;
        RECT 18.655 -23.405 18.885 -23.300 ;
        RECT 20.235 -23.405 20.465 -23.300 ;
        RECT 21.815 -23.405 22.045 -23.300 ;
        RECT 23.395 -23.405 23.625 -23.300 ;
        RECT 24.975 -23.405 25.205 -23.300 ;
        RECT 26.555 -23.405 26.785 -23.300 ;
        RECT 28.135 -23.405 28.365 -23.300 ;
        RECT 29.715 -23.405 29.945 -23.300 ;
        RECT 31.295 -23.405 31.525 -23.300 ;
        RECT 32.875 -23.405 33.105 -23.300 ;
        RECT 14.170 -23.670 18.180 -23.660 ;
        RECT 14.170 -23.960 33.970 -23.670 ;
        RECT 14.170 -24.350 15.400 -23.960 ;
        RECT 17.840 -23.970 33.970 -23.960 ;
        RECT 18.275 -24.210 33.485 -24.205 ;
        RECT 37.230 -24.210 37.530 -12.620 ;
        RECT 17.840 -24.510 37.530 -24.210 ;
      LAYER met2 ;
        RECT 11.130 0.000 163.130 107.285 ;
        RECT 16.450 -13.660 35.110 -9.850 ;
        RECT 14.190 -18.260 15.410 -16.760 ;
        RECT 16.320 -17.970 35.220 -13.660 ;
        RECT 16.340 -23.300 35.240 -18.990 ;
        RECT 16.380 -26.290 35.040 -23.300 ;
      LAYER met3 ;
        RECT 7.630 0.000 164.960 108.150 ;
        RECT 164.430 -4.855 164.940 0.000 ;
        RECT 64.610 -5.375 164.945 -4.855 ;
        RECT 16.390 -14.120 35.040 -9.860 ;
        RECT 64.680 -17.125 65.200 -5.375 ;
        RECT 14.250 -17.670 65.215 -17.125 ;
        RECT 16.390 -27.220 35.040 -22.960 ;
      LAYER met4 ;
        RECT 0.000 97.340 7.270 108.150 ;
        RECT 8.370 100.060 10.950 108.150 ;
        RECT 12.050 100.060 14.630 108.150 ;
        RECT 15.730 100.060 18.310 108.150 ;
        RECT 8.370 97.340 18.310 100.060 ;
        RECT 19.410 100.060 21.990 108.150 ;
        RECT 23.090 104.140 25.670 108.150 ;
        RECT 26.770 104.140 29.350 108.150 ;
        RECT 23.090 100.060 29.350 104.140 ;
        RECT 30.450 100.060 33.030 108.150 ;
        RECT 34.130 106.860 36.710 108.150 ;
        RECT 37.810 106.860 40.390 108.150 ;
        RECT 41.490 106.860 44.070 108.150 ;
        RECT 45.170 106.860 47.750 108.150 ;
        RECT 34.130 104.000 47.750 106.860 ;
        RECT 34.130 100.060 43.530 104.000 ;
        RECT 19.410 97.340 43.530 100.060 ;
        RECT 0.000 4.800 43.530 97.340 ;
        RECT 45.930 97.340 47.750 104.000 ;
        RECT 48.850 106.860 51.430 108.150 ;
        RECT 52.530 106.860 55.110 108.150 ;
        RECT 48.850 106.180 55.110 106.860 ;
        RECT 56.210 106.180 58.790 108.150 ;
        RECT 48.850 100.060 58.790 106.180 ;
        RECT 59.890 102.100 62.470 108.150 ;
        RECT 63.570 106.860 66.150 108.150 ;
        RECT 67.250 106.860 69.830 108.150 ;
        RECT 70.930 106.860 73.510 108.150 ;
        RECT 63.570 102.780 73.510 106.860 ;
        RECT 74.610 106.860 77.190 108.150 ;
        RECT 78.290 106.860 80.870 108.150 ;
        RECT 74.610 102.780 80.870 106.860 ;
        RECT 81.970 104.140 84.550 108.150 ;
        RECT 85.650 106.860 88.230 108.150 ;
        RECT 89.330 106.860 91.910 108.150 ;
        RECT 85.650 104.140 91.910 106.860 ;
        RECT 81.970 104.000 91.910 104.140 ;
        RECT 81.970 102.780 82.740 104.000 ;
        RECT 63.570 102.100 82.740 102.780 ;
        RECT 59.890 100.060 82.740 102.100 ;
        RECT 48.850 97.340 82.740 100.060 ;
        RECT 45.930 4.800 82.740 97.340 ;
        RECT 85.140 102.780 91.910 104.000 ;
        RECT 93.010 106.860 95.590 108.150 ;
        RECT 96.690 106.860 99.270 108.150 ;
        RECT 100.370 106.860 102.950 108.150 ;
        RECT 104.050 106.860 106.630 108.150 ;
        RECT 107.730 106.860 110.310 108.150 ;
        RECT 111.410 106.860 113.990 108.150 ;
        RECT 115.090 106.860 117.670 108.150 ;
        RECT 93.010 102.780 117.670 106.860 ;
        RECT 85.140 102.100 117.670 102.780 ;
        RECT 118.770 106.860 121.350 108.150 ;
        RECT 122.450 107.400 125.030 108.150 ;
        RECT 126.130 107.400 128.710 108.150 ;
        RECT 129.810 107.400 132.390 108.150 ;
        RECT 133.490 107.400 136.070 108.150 ;
        RECT 137.170 107.400 139.750 108.150 ;
        RECT 140.850 107.400 143.430 108.150 ;
        RECT 144.530 107.400 147.110 108.150 ;
        RECT 148.210 107.400 150.790 108.150 ;
        RECT 122.450 106.860 150.790 107.400 ;
        RECT 151.890 106.860 154.470 108.150 ;
        RECT 155.570 106.860 158.150 108.150 ;
        RECT 118.770 106.550 158.150 106.860 ;
        RECT 159.250 106.550 161.090 108.150 ;
        RECT 118.770 104.000 161.090 106.550 ;
        RECT 118.770 102.100 121.950 104.000 ;
        RECT 85.140 4.800 121.950 102.100 ;
        RECT 124.350 4.800 161.090 104.000 ;
        RECT 0.000 0.000 161.090 4.800 ;
        RECT 23.540 -0.640 161.090 0.000 ;
        RECT 21.340 -0.860 161.090 -0.640 ;
        RECT 21.340 -2.180 44.530 -0.860 ;
        RECT 21.340 -4.970 44.840 -2.180 ;
        RECT 4.020 -11.690 12.210 -7.750 ;
        RECT 38.660 -8.030 44.840 -4.970 ;
        RECT 38.660 -8.140 48.540 -8.030 ;
        RECT -0.420 -23.390 12.210 -11.690 ;
        RECT 14.850 -14.320 48.540 -8.140 ;
        RECT 39.150 -14.870 48.540 -14.320 ;
        RECT 40.970 -15.470 48.540 -14.870 ;
        RECT 15.320 -23.390 39.150 -23.220 ;
        RECT -0.420 -25.000 39.150 -23.390 ;
        RECT 4.020 -30.480 39.150 -25.000 ;
        RECT 4.020 -30.600 17.230 -30.480 ;
        RECT 4.020 -30.860 12.210 -30.600 ;
  END
END tt_um_test
END LIBRARY

