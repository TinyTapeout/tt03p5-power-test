magic
tech sky130A
magscale 1 2
timestamp 1685872562
<< viali >>
rect 23857 20553 23891 20587
rect 25605 20553 25639 20587
rect 28457 20553 28491 20587
rect 8493 20485 8527 20519
rect 13737 20485 13771 20519
rect 2145 20417 2179 20451
rect 2789 20417 2823 20451
rect 3433 20417 3467 20451
rect 4537 20417 4571 20451
rect 5181 20417 5215 20451
rect 6009 20417 6043 20451
rect 7573 20417 7607 20451
rect 7941 20417 7975 20451
rect 10241 20417 10275 20451
rect 10885 20417 10919 20451
rect 12449 20417 12483 20451
rect 13185 20417 13219 20451
rect 17877 20417 17911 20451
rect 18061 20417 18095 20451
rect 18245 20417 18279 20451
rect 18705 20417 18739 20451
rect 19717 20417 19751 20451
rect 20269 20417 20303 20451
rect 21005 20417 21039 20451
rect 22201 20417 22235 20451
rect 22385 20417 22419 20451
rect 23213 20417 23247 20451
rect 24041 20417 24075 20451
rect 24685 20417 24719 20451
rect 25789 20417 25823 20451
rect 26433 20417 26467 20451
rect 27353 20417 27387 20451
rect 27997 20417 28031 20451
rect 28641 20417 28675 20451
rect 29929 20417 29963 20451
rect 30573 20417 30607 20451
rect 19625 20349 19659 20383
rect 21465 20349 21499 20383
rect 22017 20349 22051 20383
rect 23397 20349 23431 20383
rect 10701 20281 10735 20315
rect 19809 20281 19843 20315
rect 21373 20281 21407 20315
rect 26249 20281 26283 20315
rect 29745 20281 29779 20315
rect 9597 20213 9631 20247
rect 18889 20213 18923 20247
rect 23029 20213 23063 20247
rect 24777 20213 24811 20247
rect 25145 20213 25179 20247
rect 27169 20213 27203 20247
rect 27813 20213 27847 20247
rect 30389 20213 30423 20247
rect 1593 20009 1627 20043
rect 6745 20009 6779 20043
rect 7481 20009 7515 20043
rect 8217 20009 8251 20043
rect 9505 20009 9539 20043
rect 10149 20009 10183 20043
rect 10793 20009 10827 20043
rect 12817 20009 12851 20043
rect 24593 20009 24627 20043
rect 11345 19941 11379 19975
rect 12173 19941 12207 19975
rect 20913 19941 20947 19975
rect 22293 19873 22327 19907
rect 22661 19873 22695 19907
rect 11437 19805 11471 19839
rect 11621 19805 11655 19839
rect 12357 19805 12391 19839
rect 17785 19805 17819 19839
rect 17877 19805 17911 19839
rect 17969 19805 18003 19839
rect 18153 19805 18187 19839
rect 20729 19805 20763 19839
rect 21557 19805 21591 19839
rect 21833 19805 21867 19839
rect 22477 19805 22511 19839
rect 23121 19805 23155 19839
rect 23397 19805 23431 19839
rect 24777 19805 24811 19839
rect 25237 19805 25271 19839
rect 29009 19805 29043 19839
rect 17509 19737 17543 19771
rect 19441 19737 19475 19771
rect 19625 19737 19659 19771
rect 19809 19737 19843 19771
rect 21465 19737 21499 19771
rect 23213 19669 23247 19703
rect 25421 19669 25455 19703
rect 28825 19669 28859 19703
rect 20085 19465 20119 19499
rect 22937 19465 22971 19499
rect 18337 19329 18371 19363
rect 18705 19329 18739 19363
rect 19901 19329 19935 19363
rect 20085 19329 20119 19363
rect 20729 19329 20763 19363
rect 22017 19329 22051 19363
rect 22201 19329 22235 19363
rect 23029 19329 23063 19363
rect 23213 19329 23247 19363
rect 24317 19329 24351 19363
rect 24409 19329 24443 19363
rect 24593 19329 24627 19363
rect 24685 19329 24719 19363
rect 8953 19261 8987 19295
rect 11897 19261 11931 19295
rect 24133 19261 24167 19295
rect 17509 19193 17543 19227
rect 20913 19193 20947 19227
rect 22109 19193 22143 19227
rect 15577 18921 15611 18955
rect 22753 18921 22787 18955
rect 25145 18853 25179 18887
rect 17969 18785 18003 18819
rect 16497 18717 16531 18751
rect 17049 18717 17083 18751
rect 17877 18717 17911 18751
rect 18429 18717 18463 18751
rect 22109 18717 22143 18751
rect 22293 18717 22327 18751
rect 22937 18717 22971 18751
rect 24961 18717 24995 18751
rect 22201 18649 22235 18683
rect 24593 18649 24627 18683
rect 24777 18581 24811 18615
rect 24869 18581 24903 18615
rect 23581 18377 23615 18411
rect 23673 18241 23707 18275
rect 23489 17833 23523 17867
rect 23489 17629 23523 17663
rect 23673 17629 23707 17663
rect 22293 17153 22327 17187
rect 22385 17153 22419 17187
rect 22753 17153 22787 17187
rect 23397 17153 23431 17187
rect 23857 17153 23891 17187
rect 23121 17085 23155 17119
rect 23213 16745 23247 16779
rect 23397 16541 23431 16575
rect 24593 16541 24627 16575
rect 24777 16541 24811 16575
rect 23581 16473 23615 16507
rect 24593 16405 24627 16439
rect 17785 16201 17819 16235
rect 17969 16065 18003 16099
rect 18153 15997 18187 16031
rect 18245 15997 18279 16031
rect 24409 15113 24443 15147
rect 25421 15113 25455 15147
rect 24317 14977 24351 15011
rect 24501 14977 24535 15011
rect 24961 14977 24995 15011
rect 25053 14977 25087 15011
rect 25237 14909 25271 14943
rect 20545 14569 20579 14603
rect 20177 14433 20211 14467
rect 20361 14365 20395 14399
rect 25513 14025 25547 14059
rect 24685 13957 24719 13991
rect 25697 13957 25731 13991
rect 25881 13957 25915 13991
rect 24869 13889 24903 13923
rect 25053 13889 25087 13923
rect 24409 12801 24443 12835
rect 23949 12597 23983 12631
rect 24225 12597 24259 12631
rect 21557 12393 21591 12427
rect 21925 12393 21959 12427
rect 21741 12189 21775 12223
rect 22017 12189 22051 12223
<< metal1 >>
rect 33598 21280 33714 21294
rect 21544 21274 21620 21280
rect 21544 21216 21552 21274
rect 21612 21260 21620 21274
rect 33598 21260 33614 21280
rect 21612 21226 33614 21260
rect 21612 21216 21620 21226
rect 21544 21208 21620 21216
rect 33598 21208 33614 21226
rect 33696 21208 33714 21280
rect 33598 21192 33714 21208
rect 21726 21088 21732 21140
rect 21784 21128 21790 21140
rect 24026 21128 24032 21140
rect 21784 21100 24032 21128
rect 21784 21088 21790 21100
rect 24026 21088 24032 21100
rect 24084 21088 24090 21140
rect 18414 21020 18420 21072
rect 18472 21060 18478 21072
rect 19886 21060 19892 21072
rect 18472 21032 19892 21060
rect 18472 21020 18478 21032
rect 19886 21020 19892 21032
rect 19944 21060 19950 21072
rect 24118 21060 24124 21072
rect 19944 21032 24124 21060
rect 19944 21020 19950 21032
rect 24118 21020 24124 21032
rect 24176 21020 24182 21072
rect 18230 20952 18236 21004
rect 18288 20992 18294 21004
rect 23106 20992 23112 21004
rect 18288 20964 23112 20992
rect 18288 20952 18294 20964
rect 23106 20952 23112 20964
rect 23164 20952 23170 21004
rect 19242 20884 19248 20936
rect 19300 20924 19306 20936
rect 21082 20924 21088 20936
rect 19300 20896 21088 20924
rect 19300 20884 19306 20896
rect 21082 20884 21088 20896
rect 21140 20884 21146 20936
rect 19794 20816 19800 20868
rect 19852 20856 19858 20868
rect 22462 20856 22468 20868
rect 19852 20828 22468 20856
rect 19852 20816 19858 20828
rect 22462 20816 22468 20828
rect 22520 20856 22526 20868
rect 28442 20856 28448 20868
rect 22520 20828 28448 20856
rect 22520 20816 22526 20828
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 18046 20748 18052 20800
rect 18104 20788 18110 20800
rect 22186 20788 22192 20800
rect 18104 20760 22192 20788
rect 18104 20748 18110 20760
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 1104 20698 32632 20720
rect 1104 20646 8792 20698
rect 8844 20646 8856 20698
rect 8908 20646 8920 20698
rect 8972 20646 8984 20698
rect 9036 20646 9048 20698
rect 9100 20646 16634 20698
rect 16686 20646 16698 20698
rect 16750 20646 16762 20698
rect 16814 20646 16826 20698
rect 16878 20646 16890 20698
rect 16942 20646 24476 20698
rect 24528 20646 24540 20698
rect 24592 20646 24604 20698
rect 24656 20646 24668 20698
rect 24720 20646 24732 20698
rect 24784 20646 32318 20698
rect 32370 20646 32382 20698
rect 32434 20646 32446 20698
rect 32498 20646 32510 20698
rect 32562 20646 32574 20698
rect 32626 20646 32632 20698
rect 1104 20624 32632 20646
rect 13814 20584 13820 20596
rect 8496 20556 13820 20584
rect 8496 20525 8524 20556
rect 13814 20544 13820 20556
rect 13872 20544 13878 20596
rect 22278 20584 22284 20596
rect 17972 20556 22284 20584
rect 8481 20519 8539 20525
rect 8481 20485 8493 20519
rect 8527 20485 8539 20519
rect 12526 20516 12532 20528
rect 8481 20479 8539 20485
rect 10888 20488 12532 20516
rect 2130 20408 2136 20460
rect 2188 20408 2194 20460
rect 2774 20408 2780 20460
rect 2832 20408 2838 20460
rect 3418 20408 3424 20460
rect 3476 20408 3482 20460
rect 4522 20408 4528 20460
rect 4580 20408 4586 20460
rect 5166 20408 5172 20460
rect 5224 20408 5230 20460
rect 5994 20408 6000 20460
rect 6052 20408 6058 20460
rect 7558 20408 7564 20460
rect 7616 20408 7622 20460
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20448 7987 20451
rect 10226 20448 10232 20460
rect 7975 20420 10232 20448
rect 7975 20417 7987 20420
rect 7929 20411 7987 20417
rect 10226 20408 10232 20420
rect 10284 20408 10290 20460
rect 10888 20457 10916 20488
rect 12526 20476 12532 20488
rect 12584 20516 12590 20528
rect 13725 20519 13783 20525
rect 12584 20488 13124 20516
rect 12584 20476 12590 20488
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 12434 20408 12440 20460
rect 12492 20408 12498 20460
rect 13096 20380 13124 20488
rect 13725 20485 13737 20519
rect 13771 20516 13783 20519
rect 13998 20516 14004 20528
rect 13771 20488 14004 20516
rect 13771 20485 13783 20488
rect 13725 20479 13783 20485
rect 13998 20476 14004 20488
rect 14056 20476 14062 20528
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20448 13231 20451
rect 17865 20451 17923 20457
rect 17865 20448 17877 20451
rect 13219 20420 17877 20448
rect 13219 20417 13231 20420
rect 13173 20411 13231 20417
rect 17865 20417 17877 20420
rect 17911 20417 17923 20451
rect 17865 20411 17923 20417
rect 17972 20380 18000 20556
rect 22278 20544 22284 20556
rect 22336 20544 22342 20596
rect 23750 20584 23756 20596
rect 23124 20556 23756 20584
rect 22646 20516 22652 20528
rect 18064 20488 22652 20516
rect 18064 20457 18092 20488
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18230 20408 18236 20460
rect 18288 20408 18294 20460
rect 18693 20451 18751 20457
rect 18693 20417 18705 20451
rect 18739 20448 18751 20451
rect 19518 20448 19524 20460
rect 18739 20420 19524 20448
rect 18739 20417 18751 20420
rect 18693 20411 18751 20417
rect 19518 20408 19524 20420
rect 19576 20408 19582 20460
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20448 19763 20451
rect 20162 20448 20168 20460
rect 19751 20420 20168 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20254 20408 20260 20460
rect 20312 20408 20318 20460
rect 20346 20408 20352 20460
rect 20404 20448 20410 20460
rect 22204 20457 22232 20488
rect 22646 20476 22652 20488
rect 22704 20476 22710 20528
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20404 20420 21005 20448
rect 20404 20408 20410 20420
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 22189 20451 22247 20457
rect 20993 20411 21051 20417
rect 21100 20420 22140 20448
rect 13096 20352 18000 20380
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 18196 20352 19625 20380
rect 18196 20340 18202 20352
rect 19613 20349 19625 20352
rect 19659 20380 19671 20383
rect 21100 20380 21128 20420
rect 19659 20352 21128 20380
rect 19659 20349 19671 20352
rect 19613 20343 19671 20349
rect 21174 20340 21180 20392
rect 21232 20380 21238 20392
rect 21453 20383 21511 20389
rect 21453 20380 21465 20383
rect 21232 20352 21465 20380
rect 21232 20340 21238 20352
rect 21453 20349 21465 20352
rect 21499 20349 21511 20383
rect 21453 20343 21511 20349
rect 21910 20340 21916 20392
rect 21968 20380 21974 20392
rect 22005 20383 22063 20389
rect 22005 20380 22017 20383
rect 21968 20352 22017 20380
rect 21968 20340 21974 20352
rect 22005 20349 22017 20352
rect 22051 20349 22063 20383
rect 22112 20380 22140 20420
rect 22189 20417 22201 20451
rect 22235 20417 22247 20451
rect 22189 20411 22247 20417
rect 22370 20408 22376 20460
rect 22428 20408 22434 20460
rect 22738 20380 22744 20392
rect 22112 20352 22744 20380
rect 22005 20343 22063 20349
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 10689 20315 10747 20321
rect 10689 20281 10701 20315
rect 10735 20312 10747 20315
rect 12802 20312 12808 20324
rect 10735 20284 12808 20312
rect 10735 20281 10747 20284
rect 10689 20275 10747 20281
rect 12802 20272 12808 20284
rect 12860 20272 12866 20324
rect 19797 20315 19855 20321
rect 19797 20281 19809 20315
rect 19843 20312 19855 20315
rect 19886 20312 19892 20324
rect 19843 20284 19892 20312
rect 19843 20281 19855 20284
rect 19797 20275 19855 20281
rect 19886 20272 19892 20284
rect 19944 20272 19950 20324
rect 20162 20272 20168 20324
rect 20220 20312 20226 20324
rect 20990 20312 20996 20324
rect 20220 20284 20996 20312
rect 20220 20272 20226 20284
rect 20990 20272 20996 20284
rect 21048 20272 21054 20324
rect 21361 20315 21419 20321
rect 21361 20281 21373 20315
rect 21407 20312 21419 20315
rect 23124 20312 23152 20556
rect 23750 20544 23756 20556
rect 23808 20544 23814 20596
rect 23842 20544 23848 20596
rect 23900 20544 23906 20596
rect 24302 20544 24308 20596
rect 24360 20584 24366 20596
rect 25593 20587 25651 20593
rect 25593 20584 25605 20587
rect 24360 20556 25605 20584
rect 24360 20544 24366 20556
rect 25593 20553 25605 20556
rect 25639 20553 25651 20587
rect 25593 20547 25651 20553
rect 28442 20544 28448 20596
rect 28500 20544 28506 20596
rect 23658 20476 23664 20528
rect 23716 20516 23722 20528
rect 23716 20488 25820 20516
rect 23716 20476 23722 20488
rect 23201 20451 23259 20457
rect 23201 20417 23213 20451
rect 23247 20448 23259 20451
rect 23566 20448 23572 20460
rect 23247 20420 23572 20448
rect 23247 20417 23259 20420
rect 23201 20411 23259 20417
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24210 20408 24216 20460
rect 24268 20448 24274 20460
rect 25792 20457 25820 20488
rect 24673 20451 24731 20457
rect 24673 20448 24685 20451
rect 24268 20420 24685 20448
rect 24268 20408 24274 20420
rect 24673 20417 24685 20420
rect 24719 20417 24731 20451
rect 24673 20411 24731 20417
rect 25777 20451 25835 20457
rect 25777 20417 25789 20451
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 25866 20408 25872 20460
rect 25924 20448 25930 20460
rect 26421 20451 26479 20457
rect 26421 20448 26433 20451
rect 25924 20420 26433 20448
rect 25924 20408 25930 20420
rect 26421 20417 26433 20420
rect 26467 20417 26479 20451
rect 26421 20411 26479 20417
rect 27338 20408 27344 20460
rect 27396 20408 27402 20460
rect 27430 20408 27436 20460
rect 27488 20448 27494 20460
rect 27985 20451 28043 20457
rect 27985 20448 27997 20451
rect 27488 20420 27997 20448
rect 27488 20408 27494 20420
rect 27985 20417 27997 20420
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 28626 20408 28632 20460
rect 28684 20408 28690 20460
rect 29914 20408 29920 20460
rect 29972 20408 29978 20460
rect 30282 20408 30288 20460
rect 30340 20448 30346 20460
rect 30561 20451 30619 20457
rect 30561 20448 30573 20451
rect 30340 20420 30573 20448
rect 30340 20408 30346 20420
rect 30561 20417 30573 20420
rect 30607 20417 30619 20451
rect 30561 20411 30619 20417
rect 23382 20340 23388 20392
rect 23440 20340 23446 20392
rect 24486 20340 24492 20392
rect 24544 20380 24550 20392
rect 24544 20352 29776 20380
rect 24544 20340 24550 20352
rect 21407 20284 23152 20312
rect 21407 20281 21419 20284
rect 21361 20275 21419 20281
rect 23474 20272 23480 20324
rect 23532 20312 23538 20324
rect 29748 20321 29776 20352
rect 26237 20315 26295 20321
rect 26237 20312 26249 20315
rect 23532 20284 26249 20312
rect 23532 20272 23538 20284
rect 26237 20281 26249 20284
rect 26283 20281 26295 20315
rect 26237 20275 26295 20281
rect 29733 20315 29791 20321
rect 29733 20281 29745 20315
rect 29779 20281 29791 20315
rect 29733 20275 29791 20281
rect 9585 20247 9643 20253
rect 9585 20213 9597 20247
rect 9631 20244 9643 20247
rect 11422 20244 11428 20256
rect 9631 20216 11428 20244
rect 9631 20213 9643 20216
rect 9585 20207 9643 20213
rect 11422 20204 11428 20216
rect 11480 20204 11486 20256
rect 18874 20204 18880 20256
rect 18932 20204 18938 20256
rect 20254 20204 20260 20256
rect 20312 20244 20318 20256
rect 23017 20247 23075 20253
rect 23017 20244 23029 20247
rect 20312 20216 23029 20244
rect 20312 20204 20318 20216
rect 23017 20213 23029 20216
rect 23063 20244 23075 20247
rect 24765 20247 24823 20253
rect 24765 20244 24777 20247
rect 23063 20216 24777 20244
rect 23063 20213 23075 20216
rect 23017 20207 23075 20213
rect 24765 20213 24777 20216
rect 24811 20244 24823 20247
rect 24854 20244 24860 20256
rect 24811 20216 24860 20244
rect 24811 20213 24823 20216
rect 24765 20207 24823 20213
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 25130 20204 25136 20256
rect 25188 20204 25194 20256
rect 27154 20204 27160 20256
rect 27212 20204 27218 20256
rect 27798 20204 27804 20256
rect 27856 20204 27862 20256
rect 30374 20204 30380 20256
rect 30432 20204 30438 20256
rect 1104 20154 32476 20176
rect 1104 20102 4871 20154
rect 4923 20102 4935 20154
rect 4987 20102 4999 20154
rect 5051 20102 5063 20154
rect 5115 20102 5127 20154
rect 5179 20102 12713 20154
rect 12765 20102 12777 20154
rect 12829 20102 12841 20154
rect 12893 20102 12905 20154
rect 12957 20102 12969 20154
rect 13021 20102 20555 20154
rect 20607 20102 20619 20154
rect 20671 20102 20683 20154
rect 20735 20102 20747 20154
rect 20799 20102 20811 20154
rect 20863 20102 28397 20154
rect 28449 20102 28461 20154
rect 28513 20102 28525 20154
rect 28577 20102 28589 20154
rect 28641 20102 28653 20154
rect 28705 20102 32476 20154
rect 1104 20080 32476 20102
rect 1578 20000 1584 20052
rect 1636 20000 1642 20052
rect 6730 20000 6736 20052
rect 6788 20000 6794 20052
rect 7466 20000 7472 20052
rect 7524 20000 7530 20052
rect 8202 20000 8208 20052
rect 8260 20000 8266 20052
rect 9493 20043 9551 20049
rect 9493 20009 9505 20043
rect 9539 20040 9551 20043
rect 9674 20040 9680 20052
rect 9539 20012 9680 20040
rect 9539 20009 9551 20012
rect 9493 20003 9551 20009
rect 9674 20000 9680 20012
rect 9732 20000 9738 20052
rect 10134 20000 10140 20052
rect 10192 20000 10198 20052
rect 10781 20043 10839 20049
rect 10781 20009 10793 20043
rect 10827 20040 10839 20043
rect 11054 20040 11060 20052
rect 10827 20012 11060 20040
rect 10827 20009 10839 20012
rect 10781 20003 10839 20009
rect 11054 20000 11060 20012
rect 11112 20000 11118 20052
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 12805 20043 12863 20049
rect 12805 20040 12817 20043
rect 12676 20012 12817 20040
rect 12676 20000 12682 20012
rect 12805 20009 12817 20012
rect 12851 20009 12863 20043
rect 12805 20003 12863 20009
rect 17862 20000 17868 20052
rect 17920 20040 17926 20052
rect 18414 20040 18420 20052
rect 17920 20012 18420 20040
rect 17920 20000 17926 20012
rect 18414 20000 18420 20012
rect 18472 20000 18478 20052
rect 18874 20000 18880 20052
rect 18932 20040 18938 20052
rect 18932 20012 22692 20040
rect 18932 20000 18938 20012
rect 7558 19932 7564 19984
rect 7616 19972 7622 19984
rect 11333 19975 11391 19981
rect 11333 19972 11345 19975
rect 7616 19944 11345 19972
rect 7616 19932 7622 19944
rect 11333 19941 11345 19944
rect 11379 19941 11391 19975
rect 11333 19935 11391 19941
rect 12161 19975 12219 19981
rect 12161 19941 12173 19975
rect 12207 19972 12219 19975
rect 15746 19972 15752 19984
rect 12207 19944 15752 19972
rect 12207 19941 12219 19944
rect 12161 19935 12219 19941
rect 15746 19932 15752 19944
rect 15804 19932 15810 19984
rect 20806 19972 20812 19984
rect 16960 19944 20812 19972
rect 12526 19904 12532 19916
rect 11624 19876 12532 19904
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 11624 19845 11652 19876
rect 12526 19864 12532 19876
rect 12584 19864 12590 19916
rect 11609 19839 11667 19845
rect 11609 19805 11621 19839
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 12345 19839 12403 19845
rect 12345 19805 12357 19839
rect 12391 19836 12403 19839
rect 16960 19836 16988 19944
rect 20806 19932 20812 19944
rect 20864 19932 20870 19984
rect 20901 19975 20959 19981
rect 20901 19941 20913 19975
rect 20947 19972 20959 19975
rect 21082 19972 21088 19984
rect 20947 19944 21088 19972
rect 20947 19941 20959 19944
rect 20901 19935 20959 19941
rect 21082 19932 21088 19944
rect 21140 19932 21146 19984
rect 17218 19864 17224 19916
rect 17276 19904 17282 19916
rect 17276 19876 21036 19904
rect 17276 19864 17282 19876
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 12391 19808 16988 19836
rect 17420 19808 17785 19836
rect 12391 19805 12403 19808
rect 12345 19799 12403 19805
rect 17420 19700 17448 19808
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 17957 19839 18015 19845
rect 17957 19805 17969 19839
rect 18003 19836 18015 19839
rect 18046 19836 18052 19848
rect 18003 19808 18052 19836
rect 18003 19805 18015 19808
rect 17957 19799 18015 19805
rect 18046 19796 18052 19808
rect 18104 19796 18110 19848
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19836 18199 19839
rect 19242 19836 19248 19848
rect 18187 19808 19248 19836
rect 18187 19805 18199 19808
rect 18141 19799 18199 19805
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 20346 19836 20352 19848
rect 19352 19808 20352 19836
rect 17497 19771 17555 19777
rect 17497 19737 17509 19771
rect 17543 19768 17555 19771
rect 19352 19768 19380 19808
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 20438 19796 20444 19848
rect 20496 19836 20502 19848
rect 20717 19839 20775 19845
rect 20717 19836 20729 19839
rect 20496 19808 20729 19836
rect 20496 19796 20502 19808
rect 20717 19805 20729 19808
rect 20763 19805 20775 19839
rect 21008 19836 21036 19876
rect 21192 19876 22232 19904
rect 21192 19836 21220 19876
rect 21008 19808 21220 19836
rect 20717 19799 20775 19805
rect 21542 19796 21548 19848
rect 21600 19796 21606 19848
rect 21818 19796 21824 19848
rect 21876 19796 21882 19848
rect 17543 19740 19380 19768
rect 19429 19771 19487 19777
rect 17543 19737 17555 19740
rect 17497 19731 17555 19737
rect 19429 19737 19441 19771
rect 19475 19768 19487 19771
rect 19518 19768 19524 19780
rect 19475 19740 19524 19768
rect 19475 19737 19487 19740
rect 19429 19731 19487 19737
rect 19518 19728 19524 19740
rect 19576 19728 19582 19780
rect 19613 19771 19671 19777
rect 19613 19737 19625 19771
rect 19659 19737 19671 19771
rect 19613 19731 19671 19737
rect 18046 19700 18052 19712
rect 17420 19672 18052 19700
rect 18046 19660 18052 19672
rect 18104 19660 18110 19712
rect 19628 19700 19656 19731
rect 19794 19728 19800 19780
rect 19852 19728 19858 19780
rect 19978 19728 19984 19780
rect 20036 19768 20042 19780
rect 21453 19771 21511 19777
rect 21453 19768 21465 19771
rect 20036 19740 21465 19768
rect 20036 19728 20042 19740
rect 21453 19737 21465 19740
rect 21499 19737 21511 19771
rect 22204 19768 22232 19876
rect 22278 19864 22284 19916
rect 22336 19864 22342 19916
rect 22664 19913 22692 20012
rect 23382 20000 23388 20052
rect 23440 20040 23446 20052
rect 24581 20043 24639 20049
rect 24581 20040 24593 20043
rect 23440 20012 24593 20040
rect 23440 20000 23446 20012
rect 24581 20009 24593 20012
rect 24627 20009 24639 20043
rect 24581 20003 24639 20009
rect 22830 19932 22836 19984
rect 22888 19972 22894 19984
rect 23474 19972 23480 19984
rect 22888 19944 23480 19972
rect 22888 19932 22894 19944
rect 22649 19907 22707 19913
rect 22649 19873 22661 19907
rect 22695 19904 22707 19907
rect 22695 19876 23152 19904
rect 22695 19873 22707 19876
rect 22649 19867 22707 19873
rect 22465 19839 22523 19845
rect 22465 19805 22477 19839
rect 22511 19836 22523 19839
rect 22830 19836 22836 19848
rect 22511 19808 22836 19836
rect 22511 19805 22523 19808
rect 22465 19799 22523 19805
rect 22830 19796 22836 19808
rect 22888 19796 22894 19848
rect 23124 19845 23152 19876
rect 23400 19845 23428 19944
rect 23474 19932 23480 19944
rect 23532 19932 23538 19984
rect 23934 19932 23940 19984
rect 23992 19972 23998 19984
rect 27798 19972 27804 19984
rect 23992 19944 27804 19972
rect 23992 19932 23998 19944
rect 27798 19932 27804 19944
rect 27856 19932 27862 19984
rect 24394 19864 24400 19916
rect 24452 19904 24458 19916
rect 24452 19876 25268 19904
rect 24452 19864 24458 19876
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19805 23167 19839
rect 23109 19799 23167 19805
rect 23385 19839 23443 19845
rect 23385 19805 23397 19839
rect 23431 19805 23443 19839
rect 23385 19799 23443 19805
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 25240 19845 25268 19876
rect 25225 19839 25283 19845
rect 25225 19805 25237 19839
rect 25271 19805 25283 19839
rect 25225 19799 25283 19805
rect 28810 19796 28816 19848
rect 28868 19836 28874 19848
rect 28997 19839 29055 19845
rect 28997 19836 29009 19839
rect 28868 19808 29009 19836
rect 28868 19796 28874 19808
rect 28997 19805 29009 19808
rect 29043 19805 29055 19839
rect 28997 19799 29055 19805
rect 23566 19768 23572 19780
rect 22204 19740 23244 19768
rect 21453 19731 21511 19737
rect 21634 19700 21640 19712
rect 19628 19672 21640 19700
rect 21634 19660 21640 19672
rect 21692 19660 21698 19712
rect 23216 19709 23244 19740
rect 23308 19740 23572 19768
rect 23308 19712 23336 19740
rect 23566 19728 23572 19740
rect 23624 19768 23630 19780
rect 23624 19740 28856 19768
rect 23624 19728 23630 19740
rect 23201 19703 23259 19709
rect 23201 19669 23213 19703
rect 23247 19669 23259 19703
rect 23201 19663 23259 19669
rect 23290 19660 23296 19712
rect 23348 19660 23354 19712
rect 25406 19660 25412 19712
rect 25464 19660 25470 19712
rect 28828 19709 28856 19740
rect 28813 19703 28871 19709
rect 28813 19669 28825 19703
rect 28859 19669 28871 19703
rect 28813 19663 28871 19669
rect 1104 19610 32632 19632
rect 1104 19558 8792 19610
rect 8844 19558 8856 19610
rect 8908 19558 8920 19610
rect 8972 19558 8984 19610
rect 9036 19558 9048 19610
rect 9100 19558 16634 19610
rect 16686 19558 16698 19610
rect 16750 19558 16762 19610
rect 16814 19558 16826 19610
rect 16878 19558 16890 19610
rect 16942 19558 24476 19610
rect 24528 19558 24540 19610
rect 24592 19558 24604 19610
rect 24656 19558 24668 19610
rect 24720 19558 24732 19610
rect 24784 19558 32318 19610
rect 32370 19558 32382 19610
rect 32434 19558 32446 19610
rect 32498 19558 32510 19610
rect 32562 19558 32574 19610
rect 32626 19558 32632 19610
rect 1104 19536 32632 19558
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 17218 19496 17224 19508
rect 11480 19468 17224 19496
rect 11480 19456 11486 19468
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 18046 19456 18052 19508
rect 18104 19496 18110 19508
rect 19886 19496 19892 19508
rect 18104 19468 19892 19496
rect 18104 19456 18110 19468
rect 19886 19456 19892 19468
rect 19944 19456 19950 19508
rect 20073 19499 20131 19505
rect 20073 19465 20085 19499
rect 20119 19496 20131 19499
rect 20119 19468 21772 19496
rect 20119 19465 20131 19468
rect 20073 19459 20131 19465
rect 19794 19428 19800 19440
rect 18340 19400 19800 19428
rect 18340 19369 18368 19400
rect 19794 19388 19800 19400
rect 19852 19388 19858 19440
rect 21744 19428 21772 19468
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 22094 19496 22100 19508
rect 22060 19468 22100 19496
rect 22060 19456 22066 19468
rect 22094 19456 22100 19468
rect 22152 19456 22158 19508
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 22925 19499 22983 19505
rect 22925 19496 22937 19499
rect 22796 19468 22937 19496
rect 22796 19456 22802 19468
rect 22925 19465 22937 19468
rect 22971 19465 22983 19499
rect 22925 19459 22983 19465
rect 23014 19456 23020 19508
rect 23072 19496 23078 19508
rect 27154 19496 27160 19508
rect 23072 19468 27160 19496
rect 23072 19456 23078 19468
rect 27154 19456 27160 19468
rect 27212 19456 27218 19508
rect 23290 19428 23296 19440
rect 19904 19400 21588 19428
rect 21744 19400 22968 19428
rect 19904 19369 19932 19400
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 18693 19363 18751 19369
rect 18693 19329 18705 19363
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19360 20131 19363
rect 20717 19363 20775 19369
rect 20119 19332 20668 19360
rect 20119 19329 20131 19332
rect 20073 19323 20131 19329
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19292 8999 19295
rect 9122 19292 9128 19304
rect 8987 19264 9128 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 11882 19252 11888 19304
rect 11940 19252 11946 19304
rect 18708 19292 18736 19323
rect 20640 19304 20668 19332
rect 20717 19329 20729 19363
rect 20763 19360 20775 19363
rect 20898 19360 20904 19372
rect 20763 19332 20904 19360
rect 20763 19329 20775 19332
rect 20717 19323 20775 19329
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 19978 19292 19984 19304
rect 18708 19264 19984 19292
rect 19978 19252 19984 19264
rect 20036 19252 20042 19304
rect 20622 19252 20628 19304
rect 20680 19292 20686 19304
rect 20680 19264 20944 19292
rect 20680 19252 20686 19264
rect 10226 19184 10232 19236
rect 10284 19224 10290 19236
rect 17218 19224 17224 19236
rect 10284 19196 17224 19224
rect 10284 19184 10290 19196
rect 17218 19184 17224 19196
rect 17276 19184 17282 19236
rect 17494 19184 17500 19236
rect 17552 19184 17558 19236
rect 20916 19233 20944 19264
rect 21450 19252 21456 19304
rect 21508 19292 21514 19304
rect 21560 19292 21588 19400
rect 22005 19364 22063 19369
rect 22005 19363 22140 19364
rect 22005 19329 22017 19363
rect 22051 19336 22140 19363
rect 22051 19332 22073 19336
rect 22051 19329 22063 19332
rect 22005 19323 22063 19329
rect 21508 19264 21588 19292
rect 21508 19252 21514 19264
rect 21634 19252 21640 19304
rect 21692 19292 21698 19304
rect 22112 19292 22140 19336
rect 22189 19363 22247 19369
rect 22189 19329 22201 19363
rect 22235 19360 22247 19363
rect 22462 19360 22468 19372
rect 22235 19332 22468 19360
rect 22235 19329 22247 19332
rect 22189 19323 22247 19329
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 22738 19292 22744 19304
rect 21692 19264 22744 19292
rect 21692 19252 21698 19264
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 22940 19292 22968 19400
rect 23032 19400 23296 19428
rect 23032 19369 23060 19400
rect 23290 19388 23296 19400
rect 23348 19388 23354 19440
rect 23658 19388 23664 19440
rect 23716 19428 23722 19440
rect 23716 19400 24440 19428
rect 23716 19388 23722 19400
rect 23017 19363 23075 19369
rect 23017 19329 23029 19363
rect 23063 19329 23075 19363
rect 23017 19323 23075 19329
rect 23201 19363 23259 19369
rect 23201 19329 23213 19363
rect 23247 19360 23259 19363
rect 23382 19360 23388 19372
rect 23247 19332 23388 19360
rect 23247 19329 23259 19332
rect 23201 19323 23259 19329
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 24210 19360 24216 19372
rect 23492 19332 24216 19360
rect 23290 19292 23296 19304
rect 22940 19264 23296 19292
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 23492 19292 23520 19332
rect 24210 19320 24216 19332
rect 24268 19360 24274 19372
rect 24412 19369 24440 19400
rect 24305 19363 24363 19369
rect 24305 19360 24317 19363
rect 24268 19332 24317 19360
rect 24268 19320 24274 19332
rect 24305 19329 24317 19332
rect 24351 19329 24363 19363
rect 24305 19323 24363 19329
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19329 24455 19363
rect 24581 19363 24639 19369
rect 24581 19360 24593 19363
rect 24397 19323 24455 19329
rect 24504 19332 24593 19360
rect 23400 19264 23520 19292
rect 20901 19227 20959 19233
rect 20901 19193 20913 19227
rect 20947 19193 20959 19227
rect 20901 19187 20959 19193
rect 22097 19227 22155 19233
rect 22097 19193 22109 19227
rect 22143 19224 22155 19227
rect 22186 19224 22192 19236
rect 22143 19196 22192 19224
rect 22143 19193 22155 19196
rect 22097 19187 22155 19193
rect 22186 19184 22192 19196
rect 22244 19224 22250 19236
rect 23400 19224 23428 19264
rect 23750 19252 23756 19304
rect 23808 19292 23814 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23808 19264 24133 19292
rect 23808 19252 23814 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24504 19292 24532 19332
rect 24581 19329 24593 19332
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 24673 19363 24731 19369
rect 24673 19329 24685 19363
rect 24719 19360 24731 19363
rect 24854 19360 24860 19372
rect 24719 19332 24860 19360
rect 24719 19329 24731 19332
rect 24673 19323 24731 19329
rect 24854 19320 24860 19332
rect 24912 19320 24918 19372
rect 24121 19255 24179 19261
rect 24228 19264 24532 19292
rect 24228 19236 24256 19264
rect 22244 19196 23428 19224
rect 22244 19184 22250 19196
rect 24210 19184 24216 19236
rect 24268 19184 24274 19236
rect 21450 19116 21456 19168
rect 21508 19156 21514 19168
rect 22278 19156 22284 19168
rect 21508 19128 22284 19156
rect 21508 19116 21514 19128
rect 22278 19116 22284 19128
rect 22336 19156 22342 19168
rect 23014 19156 23020 19168
rect 22336 19128 23020 19156
rect 22336 19116 22342 19128
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 1104 19066 32476 19088
rect 1104 19014 4871 19066
rect 4923 19014 4935 19066
rect 4987 19014 4999 19066
rect 5051 19014 5063 19066
rect 5115 19014 5127 19066
rect 5179 19014 12713 19066
rect 12765 19014 12777 19066
rect 12829 19014 12841 19066
rect 12893 19014 12905 19066
rect 12957 19014 12969 19066
rect 13021 19014 20555 19066
rect 20607 19014 20619 19066
rect 20671 19014 20683 19066
rect 20735 19014 20747 19066
rect 20799 19014 20811 19066
rect 20863 19014 28397 19066
rect 28449 19014 28461 19066
rect 28513 19014 28525 19066
rect 28577 19014 28589 19066
rect 28641 19014 28653 19066
rect 28705 19014 32476 19066
rect 1104 18992 32476 19014
rect 15562 18912 15568 18964
rect 15620 18912 15626 18964
rect 22738 18912 22744 18964
rect 22796 18912 22802 18964
rect 17218 18844 17224 18896
rect 17276 18884 17282 18896
rect 25133 18887 25191 18893
rect 25133 18884 25145 18887
rect 17276 18856 25145 18884
rect 17276 18844 17282 18856
rect 25133 18853 25145 18856
rect 25179 18853 25191 18887
rect 25133 18847 25191 18853
rect 17954 18776 17960 18828
rect 18012 18776 18018 18828
rect 23106 18776 23112 18828
rect 23164 18816 23170 18828
rect 23164 18788 25084 18816
rect 23164 18776 23170 18788
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18717 16543 18751
rect 16485 18711 16543 18717
rect 16500 18680 16528 18711
rect 17034 18708 17040 18760
rect 17092 18708 17098 18760
rect 17862 18708 17868 18760
rect 17920 18708 17926 18760
rect 18414 18708 18420 18760
rect 18472 18708 18478 18760
rect 22094 18708 22100 18760
rect 22152 18708 22158 18760
rect 22278 18708 22284 18760
rect 22336 18708 22342 18760
rect 22922 18708 22928 18760
rect 22980 18708 22986 18760
rect 23474 18708 23480 18760
rect 23532 18748 23538 18760
rect 23750 18748 23756 18760
rect 23532 18720 23756 18748
rect 23532 18708 23538 18720
rect 23750 18708 23756 18720
rect 23808 18748 23814 18760
rect 24949 18751 25007 18757
rect 24949 18748 24961 18751
rect 23808 18720 24961 18748
rect 23808 18708 23814 18720
rect 24949 18717 24961 18720
rect 24995 18717 25007 18751
rect 24949 18711 25007 18717
rect 21910 18680 21916 18692
rect 16500 18652 21916 18680
rect 21910 18640 21916 18652
rect 21968 18640 21974 18692
rect 22189 18683 22247 18689
rect 22189 18649 22201 18683
rect 22235 18680 22247 18683
rect 24210 18680 24216 18692
rect 22235 18652 24216 18680
rect 22235 18649 22247 18652
rect 22189 18643 22247 18649
rect 24210 18640 24216 18652
rect 24268 18680 24274 18692
rect 24581 18683 24639 18689
rect 24581 18680 24593 18683
rect 24268 18652 24593 18680
rect 24268 18640 24274 18652
rect 24581 18649 24593 18652
rect 24627 18649 24639 18683
rect 24581 18643 24639 18649
rect 23474 18572 23480 18624
rect 23532 18612 23538 18624
rect 24765 18615 24823 18621
rect 24765 18612 24777 18615
rect 23532 18584 24777 18612
rect 23532 18572 23538 18584
rect 24765 18581 24777 18584
rect 24811 18581 24823 18615
rect 24765 18575 24823 18581
rect 24857 18615 24915 18621
rect 24857 18581 24869 18615
rect 24903 18612 24915 18615
rect 25056 18612 25084 18788
rect 24903 18584 25084 18612
rect 24903 18581 24915 18584
rect 24857 18575 24915 18581
rect 1104 18522 32632 18544
rect 1104 18470 8792 18522
rect 8844 18470 8856 18522
rect 8908 18470 8920 18522
rect 8972 18470 8984 18522
rect 9036 18470 9048 18522
rect 9100 18470 16634 18522
rect 16686 18470 16698 18522
rect 16750 18470 16762 18522
rect 16814 18470 16826 18522
rect 16878 18470 16890 18522
rect 16942 18470 24476 18522
rect 24528 18470 24540 18522
rect 24592 18470 24604 18522
rect 24656 18470 24668 18522
rect 24720 18470 24732 18522
rect 24784 18470 32318 18522
rect 32370 18470 32382 18522
rect 32434 18470 32446 18522
rect 32498 18470 32510 18522
rect 32562 18470 32574 18522
rect 32626 18470 32632 18522
rect 1104 18448 32632 18470
rect 23566 18368 23572 18420
rect 23624 18368 23630 18420
rect 17034 18300 17040 18352
rect 17092 18340 17098 18352
rect 25314 18340 25320 18352
rect 17092 18312 25320 18340
rect 17092 18300 17098 18312
rect 25314 18300 25320 18312
rect 25372 18300 25378 18352
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18272 23719 18275
rect 24026 18272 24032 18284
rect 23707 18244 24032 18272
rect 23707 18241 23719 18244
rect 23661 18235 23719 18241
rect 24026 18232 24032 18244
rect 24084 18232 24090 18284
rect 1104 17978 32476 18000
rect 1104 17926 4871 17978
rect 4923 17926 4935 17978
rect 4987 17926 4999 17978
rect 5051 17926 5063 17978
rect 5115 17926 5127 17978
rect 5179 17926 12713 17978
rect 12765 17926 12777 17978
rect 12829 17926 12841 17978
rect 12893 17926 12905 17978
rect 12957 17926 12969 17978
rect 13021 17926 20555 17978
rect 20607 17926 20619 17978
rect 20671 17926 20683 17978
rect 20735 17926 20747 17978
rect 20799 17926 20811 17978
rect 20863 17926 28397 17978
rect 28449 17926 28461 17978
rect 28513 17926 28525 17978
rect 28577 17926 28589 17978
rect 28641 17926 28653 17978
rect 28705 17926 32476 17978
rect 1104 17904 32476 17926
rect 22646 17824 22652 17876
rect 22704 17864 22710 17876
rect 23474 17864 23480 17876
rect 22704 17836 23480 17864
rect 22704 17824 22710 17836
rect 23474 17824 23480 17836
rect 23532 17824 23538 17876
rect 23566 17728 23572 17740
rect 23492 17700 23572 17728
rect 23492 17669 23520 17700
rect 23566 17688 23572 17700
rect 23624 17728 23630 17740
rect 23934 17728 23940 17740
rect 23624 17700 23940 17728
rect 23624 17688 23630 17700
rect 23934 17688 23940 17700
rect 23992 17688 23998 17740
rect 23477 17663 23535 17669
rect 23477 17629 23489 17663
rect 23523 17629 23535 17663
rect 23477 17623 23535 17629
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17660 23719 17663
rect 23842 17660 23848 17672
rect 23707 17632 23848 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 1104 17434 32632 17456
rect 1104 17382 8792 17434
rect 8844 17382 8856 17434
rect 8908 17382 8920 17434
rect 8972 17382 8984 17434
rect 9036 17382 9048 17434
rect 9100 17382 16634 17434
rect 16686 17382 16698 17434
rect 16750 17382 16762 17434
rect 16814 17382 16826 17434
rect 16878 17382 16890 17434
rect 16942 17382 24476 17434
rect 24528 17382 24540 17434
rect 24592 17382 24604 17434
rect 24656 17382 24668 17434
rect 24720 17382 24732 17434
rect 24784 17382 32318 17434
rect 32370 17382 32382 17434
rect 32434 17382 32446 17434
rect 32498 17382 32510 17434
rect 32562 17382 32574 17434
rect 32626 17382 32632 17434
rect 1104 17360 32632 17382
rect 23658 17320 23664 17332
rect 22388 17292 23664 17320
rect 22388 17252 22416 17292
rect 23658 17280 23664 17292
rect 23716 17280 23722 17332
rect 25130 17252 25136 17264
rect 22296 17224 22416 17252
rect 23400 17224 25136 17252
rect 19518 17144 19524 17196
rect 19576 17184 19582 17196
rect 22296 17193 22324 17224
rect 22281 17187 22339 17193
rect 22281 17184 22293 17187
rect 19576 17156 22293 17184
rect 19576 17144 19582 17156
rect 22281 17153 22293 17156
rect 22327 17153 22339 17187
rect 22281 17147 22339 17153
rect 22370 17144 22376 17196
rect 22428 17144 22434 17196
rect 22646 17144 22652 17196
rect 22704 17184 22710 17196
rect 23400 17193 23428 17224
rect 25130 17212 25136 17224
rect 25188 17212 25194 17264
rect 22741 17187 22799 17193
rect 22741 17184 22753 17187
rect 22704 17156 22753 17184
rect 22704 17144 22710 17156
rect 22741 17153 22753 17156
rect 22787 17153 22799 17187
rect 22741 17147 22799 17153
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17153 23443 17187
rect 23385 17147 23443 17153
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17184 23903 17187
rect 23934 17184 23940 17196
rect 23891 17156 23940 17184
rect 23891 17153 23903 17156
rect 23845 17147 23903 17153
rect 23934 17144 23940 17156
rect 23992 17184 23998 17196
rect 24118 17184 24124 17196
rect 23992 17156 24124 17184
rect 23992 17144 23998 17156
rect 24118 17144 24124 17156
rect 24176 17144 24182 17196
rect 23106 17076 23112 17128
rect 23164 17076 23170 17128
rect 1104 16890 32476 16912
rect 1104 16838 4871 16890
rect 4923 16838 4935 16890
rect 4987 16838 4999 16890
rect 5051 16838 5063 16890
rect 5115 16838 5127 16890
rect 5179 16838 12713 16890
rect 12765 16838 12777 16890
rect 12829 16838 12841 16890
rect 12893 16838 12905 16890
rect 12957 16838 12969 16890
rect 13021 16838 20555 16890
rect 20607 16838 20619 16890
rect 20671 16838 20683 16890
rect 20735 16838 20747 16890
rect 20799 16838 20811 16890
rect 20863 16838 28397 16890
rect 28449 16838 28461 16890
rect 28513 16838 28525 16890
rect 28577 16838 28589 16890
rect 28641 16838 28653 16890
rect 28705 16838 32476 16890
rect 1104 16816 32476 16838
rect 22370 16736 22376 16788
rect 22428 16776 22434 16788
rect 23201 16779 23259 16785
rect 23201 16776 23213 16779
rect 22428 16748 23213 16776
rect 22428 16736 22434 16748
rect 23201 16745 23213 16748
rect 23247 16745 23259 16779
rect 23201 16739 23259 16745
rect 24302 16600 24308 16652
rect 24360 16640 24366 16652
rect 24360 16612 24624 16640
rect 24360 16600 24366 16612
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23842 16572 23848 16584
rect 23431 16544 23848 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 24596 16581 24624 16612
rect 24581 16575 24639 16581
rect 24581 16541 24593 16575
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24765 16575 24823 16581
rect 24765 16541 24777 16575
rect 24811 16541 24823 16575
rect 24765 16535 24823 16541
rect 23566 16464 23572 16516
rect 23624 16464 23630 16516
rect 24118 16464 24124 16516
rect 24176 16504 24182 16516
rect 24394 16504 24400 16516
rect 24176 16476 24400 16504
rect 24176 16464 24182 16476
rect 24394 16464 24400 16476
rect 24452 16504 24458 16516
rect 24780 16504 24808 16535
rect 24452 16476 24808 16504
rect 24452 16464 24458 16476
rect 24026 16396 24032 16448
rect 24084 16436 24090 16448
rect 24581 16439 24639 16445
rect 24581 16436 24593 16439
rect 24084 16408 24593 16436
rect 24084 16396 24090 16408
rect 24581 16405 24593 16408
rect 24627 16405 24639 16439
rect 24581 16399 24639 16405
rect 1104 16346 32632 16368
rect 1104 16294 8792 16346
rect 8844 16294 8856 16346
rect 8908 16294 8920 16346
rect 8972 16294 8984 16346
rect 9036 16294 9048 16346
rect 9100 16294 16634 16346
rect 16686 16294 16698 16346
rect 16750 16294 16762 16346
rect 16814 16294 16826 16346
rect 16878 16294 16890 16346
rect 16942 16294 24476 16346
rect 24528 16294 24540 16346
rect 24592 16294 24604 16346
rect 24656 16294 24668 16346
rect 24720 16294 24732 16346
rect 24784 16294 32318 16346
rect 32370 16294 32382 16346
rect 32434 16294 32446 16346
rect 32498 16294 32510 16346
rect 32562 16294 32574 16346
rect 32626 16294 32632 16346
rect 1104 16272 32632 16294
rect 17773 16235 17831 16241
rect 17773 16201 17785 16235
rect 17819 16232 17831 16235
rect 17862 16232 17868 16244
rect 17819 16204 17868 16232
rect 17819 16201 17831 16204
rect 17773 16195 17831 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 17957 16099 18015 16105
rect 17957 16065 17969 16099
rect 18003 16096 18015 16099
rect 20990 16096 20996 16108
rect 18003 16068 20996 16096
rect 18003 16065 18015 16068
rect 17957 16059 18015 16065
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 18138 15988 18144 16040
rect 18196 15988 18202 16040
rect 18233 16031 18291 16037
rect 18233 15997 18245 16031
rect 18279 15997 18291 16031
rect 18233 15991 18291 15997
rect 18046 15920 18052 15972
rect 18104 15960 18110 15972
rect 18248 15960 18276 15991
rect 18104 15932 18276 15960
rect 18104 15920 18110 15932
rect 1104 15802 32476 15824
rect 1104 15750 4871 15802
rect 4923 15750 4935 15802
rect 4987 15750 4999 15802
rect 5051 15750 5063 15802
rect 5115 15750 5127 15802
rect 5179 15750 12713 15802
rect 12765 15750 12777 15802
rect 12829 15750 12841 15802
rect 12893 15750 12905 15802
rect 12957 15750 12969 15802
rect 13021 15750 20555 15802
rect 20607 15750 20619 15802
rect 20671 15750 20683 15802
rect 20735 15750 20747 15802
rect 20799 15750 20811 15802
rect 20863 15750 28397 15802
rect 28449 15750 28461 15802
rect 28513 15750 28525 15802
rect 28577 15750 28589 15802
rect 28641 15750 28653 15802
rect 28705 15750 32476 15802
rect 1104 15728 32476 15750
rect 1104 15258 32632 15280
rect 1104 15206 8792 15258
rect 8844 15206 8856 15258
rect 8908 15206 8920 15258
rect 8972 15206 8984 15258
rect 9036 15206 9048 15258
rect 9100 15206 16634 15258
rect 16686 15206 16698 15258
rect 16750 15206 16762 15258
rect 16814 15206 16826 15258
rect 16878 15206 16890 15258
rect 16942 15206 24476 15258
rect 24528 15206 24540 15258
rect 24592 15206 24604 15258
rect 24656 15206 24668 15258
rect 24720 15206 24732 15258
rect 24784 15206 32318 15258
rect 32370 15206 32382 15258
rect 32434 15206 32446 15258
rect 32498 15206 32510 15258
rect 32562 15206 32574 15258
rect 32626 15206 32632 15258
rect 1104 15184 32632 15206
rect 21542 15104 21548 15156
rect 21600 15144 21606 15156
rect 24397 15147 24455 15153
rect 24397 15144 24409 15147
rect 21600 15116 24409 15144
rect 21600 15104 21606 15116
rect 24397 15113 24409 15116
rect 24443 15113 24455 15147
rect 24397 15107 24455 15113
rect 25314 15104 25320 15156
rect 25372 15144 25378 15156
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 25372 15116 25421 15144
rect 25372 15104 25378 15116
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 25409 15107 25467 15113
rect 23934 15036 23940 15088
rect 23992 15076 23998 15088
rect 23992 15048 24992 15076
rect 23992 15036 23998 15048
rect 24118 14968 24124 15020
rect 24176 15008 24182 15020
rect 24305 15011 24363 15017
rect 24305 15008 24317 15011
rect 24176 14980 24317 15008
rect 24176 14968 24182 14980
rect 24305 14977 24317 14980
rect 24351 14977 24363 15011
rect 24305 14971 24363 14977
rect 24394 14968 24400 15020
rect 24452 15008 24458 15020
rect 24964 15017 24992 15048
rect 24489 15011 24547 15017
rect 24489 15008 24501 15011
rect 24452 14980 24501 15008
rect 24452 14968 24458 14980
rect 24489 14977 24501 14980
rect 24535 14977 24547 15011
rect 24489 14971 24547 14977
rect 24949 15011 25007 15017
rect 24949 14977 24961 15011
rect 24995 14977 25007 15011
rect 24949 14971 25007 14977
rect 25041 15011 25099 15017
rect 25041 14977 25053 15011
rect 25087 15008 25099 15011
rect 25130 15008 25136 15020
rect 25087 14980 25136 15008
rect 25087 14977 25099 14980
rect 25041 14971 25099 14977
rect 25130 14968 25136 14980
rect 25188 14968 25194 15020
rect 23658 14900 23664 14952
rect 23716 14940 23722 14952
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 23716 14912 25237 14940
rect 23716 14900 23722 14912
rect 25225 14909 25237 14912
rect 25271 14909 25283 14943
rect 25225 14903 25283 14909
rect 1104 14714 32476 14736
rect 1104 14662 4871 14714
rect 4923 14662 4935 14714
rect 4987 14662 4999 14714
rect 5051 14662 5063 14714
rect 5115 14662 5127 14714
rect 5179 14662 12713 14714
rect 12765 14662 12777 14714
rect 12829 14662 12841 14714
rect 12893 14662 12905 14714
rect 12957 14662 12969 14714
rect 13021 14662 20555 14714
rect 20607 14662 20619 14714
rect 20671 14662 20683 14714
rect 20735 14662 20747 14714
rect 20799 14662 20811 14714
rect 20863 14662 28397 14714
rect 28449 14662 28461 14714
rect 28513 14662 28525 14714
rect 28577 14662 28589 14714
rect 28641 14662 28653 14714
rect 28705 14662 32476 14714
rect 1104 14640 32476 14662
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 20496 14572 20545 14600
rect 20496 14560 20502 14572
rect 20533 14569 20545 14572
rect 20579 14569 20591 14603
rect 20533 14563 20591 14569
rect 19794 14424 19800 14476
rect 19852 14464 19858 14476
rect 20162 14464 20168 14476
rect 19852 14436 20168 14464
rect 19852 14424 19858 14436
rect 20162 14424 20168 14436
rect 20220 14424 20226 14476
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14396 20407 14399
rect 25498 14396 25504 14408
rect 20395 14368 25504 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 25498 14356 25504 14368
rect 25556 14356 25562 14408
rect 1104 14170 32632 14192
rect 1104 14118 8792 14170
rect 8844 14118 8856 14170
rect 8908 14118 8920 14170
rect 8972 14118 8984 14170
rect 9036 14118 9048 14170
rect 9100 14118 16634 14170
rect 16686 14118 16698 14170
rect 16750 14118 16762 14170
rect 16814 14118 16826 14170
rect 16878 14118 16890 14170
rect 16942 14118 24476 14170
rect 24528 14118 24540 14170
rect 24592 14118 24604 14170
rect 24656 14118 24668 14170
rect 24720 14118 24732 14170
rect 24784 14118 32318 14170
rect 32370 14118 32382 14170
rect 32434 14118 32446 14170
rect 32498 14118 32510 14170
rect 32562 14118 32574 14170
rect 32626 14118 32632 14170
rect 1104 14096 32632 14118
rect 25498 14016 25504 14068
rect 25556 14016 25562 14068
rect 20162 13948 20168 14000
rect 20220 13988 20226 14000
rect 24673 13991 24731 13997
rect 24673 13988 24685 13991
rect 20220 13960 24685 13988
rect 20220 13948 20226 13960
rect 24673 13957 24685 13960
rect 24719 13957 24731 13991
rect 25406 13988 25412 14000
rect 24673 13951 24731 13957
rect 24872 13960 25412 13988
rect 24872 13929 24900 13960
rect 25406 13948 25412 13960
rect 25464 13988 25470 14000
rect 25685 13991 25743 13997
rect 25685 13988 25697 13991
rect 25464 13960 25697 13988
rect 25464 13948 25470 13960
rect 25685 13957 25697 13960
rect 25731 13957 25743 13991
rect 25685 13951 25743 13957
rect 25869 13991 25927 13997
rect 25869 13957 25881 13991
rect 25915 13988 25927 13991
rect 30374 13988 30380 14000
rect 25915 13960 30380 13988
rect 25915 13957 25927 13960
rect 25869 13951 25927 13957
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25041 13923 25099 13929
rect 25041 13889 25053 13923
rect 25087 13920 25099 13923
rect 25884 13920 25912 13951
rect 30374 13948 30380 13960
rect 30432 13948 30438 14000
rect 25087 13892 25912 13920
rect 25087 13889 25099 13892
rect 25041 13883 25099 13889
rect 1104 13626 32476 13648
rect 1104 13574 4871 13626
rect 4923 13574 4935 13626
rect 4987 13574 4999 13626
rect 5051 13574 5063 13626
rect 5115 13574 5127 13626
rect 5179 13574 12713 13626
rect 12765 13574 12777 13626
rect 12829 13574 12841 13626
rect 12893 13574 12905 13626
rect 12957 13574 12969 13626
rect 13021 13574 20555 13626
rect 20607 13574 20619 13626
rect 20671 13574 20683 13626
rect 20735 13574 20747 13626
rect 20799 13574 20811 13626
rect 20863 13574 28397 13626
rect 28449 13574 28461 13626
rect 28513 13574 28525 13626
rect 28577 13574 28589 13626
rect 28641 13574 28653 13626
rect 28705 13574 32476 13626
rect 1104 13552 32476 13574
rect 1104 13082 32632 13104
rect 1104 13030 8792 13082
rect 8844 13030 8856 13082
rect 8908 13030 8920 13082
rect 8972 13030 8984 13082
rect 9036 13030 9048 13082
rect 9100 13030 16634 13082
rect 16686 13030 16698 13082
rect 16750 13030 16762 13082
rect 16814 13030 16826 13082
rect 16878 13030 16890 13082
rect 16942 13030 24476 13082
rect 24528 13030 24540 13082
rect 24592 13030 24604 13082
rect 24656 13030 24668 13082
rect 24720 13030 24732 13082
rect 24784 13030 32318 13082
rect 32370 13030 32382 13082
rect 32434 13030 32446 13082
rect 32498 13030 32510 13082
rect 32562 13030 32574 13082
rect 32626 13030 32632 13082
rect 1104 13008 32632 13030
rect 23750 12792 23756 12844
rect 23808 12832 23814 12844
rect 24397 12835 24455 12841
rect 24397 12832 24409 12835
rect 23808 12804 24409 12832
rect 23808 12792 23814 12804
rect 24397 12801 24409 12804
rect 24443 12801 24455 12835
rect 24397 12795 24455 12801
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 23937 12631 23995 12637
rect 23937 12628 23949 12631
rect 12492 12600 23949 12628
rect 12492 12588 12498 12600
rect 23937 12597 23949 12600
rect 23983 12597 23995 12631
rect 23937 12591 23995 12597
rect 24210 12588 24216 12640
rect 24268 12588 24274 12640
rect 1104 12538 32476 12560
rect 1104 12486 4871 12538
rect 4923 12486 4935 12538
rect 4987 12486 4999 12538
rect 5051 12486 5063 12538
rect 5115 12486 5127 12538
rect 5179 12486 12713 12538
rect 12765 12486 12777 12538
rect 12829 12486 12841 12538
rect 12893 12486 12905 12538
rect 12957 12486 12969 12538
rect 13021 12486 20555 12538
rect 20607 12486 20619 12538
rect 20671 12486 20683 12538
rect 20735 12486 20747 12538
rect 20799 12486 20811 12538
rect 20863 12486 28397 12538
rect 28449 12486 28461 12538
rect 28513 12486 28525 12538
rect 28577 12486 28589 12538
rect 28641 12486 28653 12538
rect 28705 12486 32476 12538
rect 1104 12464 32476 12486
rect 20990 12384 20996 12436
rect 21048 12424 21054 12436
rect 21545 12427 21603 12433
rect 21545 12424 21557 12427
rect 21048 12396 21557 12424
rect 21048 12384 21054 12396
rect 21545 12393 21557 12396
rect 21591 12393 21603 12427
rect 21545 12387 21603 12393
rect 21634 12384 21640 12436
rect 21692 12424 21698 12436
rect 21913 12427 21971 12433
rect 21913 12424 21925 12427
rect 21692 12396 21925 12424
rect 21692 12384 21698 12396
rect 21913 12393 21925 12396
rect 21959 12393 21971 12427
rect 21913 12387 21971 12393
rect 24026 12288 24032 12300
rect 21744 12260 24032 12288
rect 21744 12229 21772 12260
rect 24026 12248 24032 12260
rect 24084 12248 24090 12300
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 22005 12223 22063 12229
rect 22005 12189 22017 12223
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 20162 12112 20168 12164
rect 20220 12152 20226 12164
rect 22020 12152 22048 12183
rect 20220 12124 22048 12152
rect 20220 12112 20226 12124
rect 1104 11994 32632 12016
rect 1104 11942 8792 11994
rect 8844 11942 8856 11994
rect 8908 11942 8920 11994
rect 8972 11942 8984 11994
rect 9036 11942 9048 11994
rect 9100 11942 16634 11994
rect 16686 11942 16698 11994
rect 16750 11942 16762 11994
rect 16814 11942 16826 11994
rect 16878 11942 16890 11994
rect 16942 11942 24476 11994
rect 24528 11942 24540 11994
rect 24592 11942 24604 11994
rect 24656 11942 24668 11994
rect 24720 11942 24732 11994
rect 24784 11942 32318 11994
rect 32370 11942 32382 11994
rect 32434 11942 32446 11994
rect 32498 11942 32510 11994
rect 32562 11942 32574 11994
rect 32626 11942 32632 11994
rect 1104 11920 32632 11942
rect 1104 11450 32476 11472
rect 1104 11398 4871 11450
rect 4923 11398 4935 11450
rect 4987 11398 4999 11450
rect 5051 11398 5063 11450
rect 5115 11398 5127 11450
rect 5179 11398 12713 11450
rect 12765 11398 12777 11450
rect 12829 11398 12841 11450
rect 12893 11398 12905 11450
rect 12957 11398 12969 11450
rect 13021 11398 20555 11450
rect 20607 11398 20619 11450
rect 20671 11398 20683 11450
rect 20735 11398 20747 11450
rect 20799 11398 20811 11450
rect 20863 11398 28397 11450
rect 28449 11398 28461 11450
rect 28513 11398 28525 11450
rect 28577 11398 28589 11450
rect 28641 11398 28653 11450
rect 28705 11398 32476 11450
rect 1104 11376 32476 11398
rect 1104 10906 32632 10928
rect 1104 10854 8792 10906
rect 8844 10854 8856 10906
rect 8908 10854 8920 10906
rect 8972 10854 8984 10906
rect 9036 10854 9048 10906
rect 9100 10854 16634 10906
rect 16686 10854 16698 10906
rect 16750 10854 16762 10906
rect 16814 10854 16826 10906
rect 16878 10854 16890 10906
rect 16942 10854 24476 10906
rect 24528 10854 24540 10906
rect 24592 10854 24604 10906
rect 24656 10854 24668 10906
rect 24720 10854 24732 10906
rect 24784 10854 32318 10906
rect 32370 10854 32382 10906
rect 32434 10854 32446 10906
rect 32498 10854 32510 10906
rect 32562 10854 32574 10906
rect 32626 10854 32632 10906
rect 1104 10832 32632 10854
rect 1104 10362 32476 10384
rect 1104 10310 4871 10362
rect 4923 10310 4935 10362
rect 4987 10310 4999 10362
rect 5051 10310 5063 10362
rect 5115 10310 5127 10362
rect 5179 10310 12713 10362
rect 12765 10310 12777 10362
rect 12829 10310 12841 10362
rect 12893 10310 12905 10362
rect 12957 10310 12969 10362
rect 13021 10310 20555 10362
rect 20607 10310 20619 10362
rect 20671 10310 20683 10362
rect 20735 10310 20747 10362
rect 20799 10310 20811 10362
rect 20863 10310 28397 10362
rect 28449 10310 28461 10362
rect 28513 10310 28525 10362
rect 28577 10310 28589 10362
rect 28641 10310 28653 10362
rect 28705 10310 32476 10362
rect 1104 10288 32476 10310
rect 1104 9818 32632 9840
rect 1104 9766 8792 9818
rect 8844 9766 8856 9818
rect 8908 9766 8920 9818
rect 8972 9766 8984 9818
rect 9036 9766 9048 9818
rect 9100 9766 16634 9818
rect 16686 9766 16698 9818
rect 16750 9766 16762 9818
rect 16814 9766 16826 9818
rect 16878 9766 16890 9818
rect 16942 9766 24476 9818
rect 24528 9766 24540 9818
rect 24592 9766 24604 9818
rect 24656 9766 24668 9818
rect 24720 9766 24732 9818
rect 24784 9766 32318 9818
rect 32370 9766 32382 9818
rect 32434 9766 32446 9818
rect 32498 9766 32510 9818
rect 32562 9766 32574 9818
rect 32626 9766 32632 9818
rect 1104 9744 32632 9766
rect 1104 9274 32476 9296
rect 1104 9222 4871 9274
rect 4923 9222 4935 9274
rect 4987 9222 4999 9274
rect 5051 9222 5063 9274
rect 5115 9222 5127 9274
rect 5179 9222 12713 9274
rect 12765 9222 12777 9274
rect 12829 9222 12841 9274
rect 12893 9222 12905 9274
rect 12957 9222 12969 9274
rect 13021 9222 20555 9274
rect 20607 9222 20619 9274
rect 20671 9222 20683 9274
rect 20735 9222 20747 9274
rect 20799 9222 20811 9274
rect 20863 9222 28397 9274
rect 28449 9222 28461 9274
rect 28513 9222 28525 9274
rect 28577 9222 28589 9274
rect 28641 9222 28653 9274
rect 28705 9222 32476 9274
rect 1104 9200 32476 9222
rect 1104 8730 32632 8752
rect 1104 8678 8792 8730
rect 8844 8678 8856 8730
rect 8908 8678 8920 8730
rect 8972 8678 8984 8730
rect 9036 8678 9048 8730
rect 9100 8678 16634 8730
rect 16686 8678 16698 8730
rect 16750 8678 16762 8730
rect 16814 8678 16826 8730
rect 16878 8678 16890 8730
rect 16942 8678 24476 8730
rect 24528 8678 24540 8730
rect 24592 8678 24604 8730
rect 24656 8678 24668 8730
rect 24720 8678 24732 8730
rect 24784 8678 32318 8730
rect 32370 8678 32382 8730
rect 32434 8678 32446 8730
rect 32498 8678 32510 8730
rect 32562 8678 32574 8730
rect 32626 8678 32632 8730
rect 1104 8656 32632 8678
rect 1104 8186 32476 8208
rect 1104 8134 4871 8186
rect 4923 8134 4935 8186
rect 4987 8134 4999 8186
rect 5051 8134 5063 8186
rect 5115 8134 5127 8186
rect 5179 8134 12713 8186
rect 12765 8134 12777 8186
rect 12829 8134 12841 8186
rect 12893 8134 12905 8186
rect 12957 8134 12969 8186
rect 13021 8134 20555 8186
rect 20607 8134 20619 8186
rect 20671 8134 20683 8186
rect 20735 8134 20747 8186
rect 20799 8134 20811 8186
rect 20863 8134 28397 8186
rect 28449 8134 28461 8186
rect 28513 8134 28525 8186
rect 28577 8134 28589 8186
rect 28641 8134 28653 8186
rect 28705 8134 32476 8186
rect 1104 8112 32476 8134
rect 1104 7642 32632 7664
rect 1104 7590 8792 7642
rect 8844 7590 8856 7642
rect 8908 7590 8920 7642
rect 8972 7590 8984 7642
rect 9036 7590 9048 7642
rect 9100 7590 16634 7642
rect 16686 7590 16698 7642
rect 16750 7590 16762 7642
rect 16814 7590 16826 7642
rect 16878 7590 16890 7642
rect 16942 7590 24476 7642
rect 24528 7590 24540 7642
rect 24592 7590 24604 7642
rect 24656 7590 24668 7642
rect 24720 7590 24732 7642
rect 24784 7590 32318 7642
rect 32370 7590 32382 7642
rect 32434 7590 32446 7642
rect 32498 7590 32510 7642
rect 32562 7590 32574 7642
rect 32626 7590 32632 7642
rect 1104 7568 32632 7590
rect 1104 7098 32476 7120
rect 1104 7046 4871 7098
rect 4923 7046 4935 7098
rect 4987 7046 4999 7098
rect 5051 7046 5063 7098
rect 5115 7046 5127 7098
rect 5179 7046 12713 7098
rect 12765 7046 12777 7098
rect 12829 7046 12841 7098
rect 12893 7046 12905 7098
rect 12957 7046 12969 7098
rect 13021 7046 20555 7098
rect 20607 7046 20619 7098
rect 20671 7046 20683 7098
rect 20735 7046 20747 7098
rect 20799 7046 20811 7098
rect 20863 7046 28397 7098
rect 28449 7046 28461 7098
rect 28513 7046 28525 7098
rect 28577 7046 28589 7098
rect 28641 7046 28653 7098
rect 28705 7046 32476 7098
rect 1104 7024 32476 7046
rect 1104 6554 32632 6576
rect 1104 6502 8792 6554
rect 8844 6502 8856 6554
rect 8908 6502 8920 6554
rect 8972 6502 8984 6554
rect 9036 6502 9048 6554
rect 9100 6502 16634 6554
rect 16686 6502 16698 6554
rect 16750 6502 16762 6554
rect 16814 6502 16826 6554
rect 16878 6502 16890 6554
rect 16942 6502 24476 6554
rect 24528 6502 24540 6554
rect 24592 6502 24604 6554
rect 24656 6502 24668 6554
rect 24720 6502 24732 6554
rect 24784 6502 32318 6554
rect 32370 6502 32382 6554
rect 32434 6502 32446 6554
rect 32498 6502 32510 6554
rect 32562 6502 32574 6554
rect 32626 6502 32632 6554
rect 1104 6480 32632 6502
rect 1104 6010 32476 6032
rect 1104 5958 4871 6010
rect 4923 5958 4935 6010
rect 4987 5958 4999 6010
rect 5051 5958 5063 6010
rect 5115 5958 5127 6010
rect 5179 5958 12713 6010
rect 12765 5958 12777 6010
rect 12829 5958 12841 6010
rect 12893 5958 12905 6010
rect 12957 5958 12969 6010
rect 13021 5958 20555 6010
rect 20607 5958 20619 6010
rect 20671 5958 20683 6010
rect 20735 5958 20747 6010
rect 20799 5958 20811 6010
rect 20863 5958 28397 6010
rect 28449 5958 28461 6010
rect 28513 5958 28525 6010
rect 28577 5958 28589 6010
rect 28641 5958 28653 6010
rect 28705 5958 32476 6010
rect 1104 5936 32476 5958
rect 1104 5466 32632 5488
rect 1104 5414 8792 5466
rect 8844 5414 8856 5466
rect 8908 5414 8920 5466
rect 8972 5414 8984 5466
rect 9036 5414 9048 5466
rect 9100 5414 16634 5466
rect 16686 5414 16698 5466
rect 16750 5414 16762 5466
rect 16814 5414 16826 5466
rect 16878 5414 16890 5466
rect 16942 5414 24476 5466
rect 24528 5414 24540 5466
rect 24592 5414 24604 5466
rect 24656 5414 24668 5466
rect 24720 5414 24732 5466
rect 24784 5414 32318 5466
rect 32370 5414 32382 5466
rect 32434 5414 32446 5466
rect 32498 5414 32510 5466
rect 32562 5414 32574 5466
rect 32626 5414 32632 5466
rect 1104 5392 32632 5414
rect 1104 4922 32476 4944
rect 1104 4870 4871 4922
rect 4923 4870 4935 4922
rect 4987 4870 4999 4922
rect 5051 4870 5063 4922
rect 5115 4870 5127 4922
rect 5179 4870 12713 4922
rect 12765 4870 12777 4922
rect 12829 4870 12841 4922
rect 12893 4870 12905 4922
rect 12957 4870 12969 4922
rect 13021 4870 20555 4922
rect 20607 4870 20619 4922
rect 20671 4870 20683 4922
rect 20735 4870 20747 4922
rect 20799 4870 20811 4922
rect 20863 4870 28397 4922
rect 28449 4870 28461 4922
rect 28513 4870 28525 4922
rect 28577 4870 28589 4922
rect 28641 4870 28653 4922
rect 28705 4870 32476 4922
rect 1104 4848 32476 4870
rect 1104 4378 32632 4400
rect 1104 4326 8792 4378
rect 8844 4326 8856 4378
rect 8908 4326 8920 4378
rect 8972 4326 8984 4378
rect 9036 4326 9048 4378
rect 9100 4326 16634 4378
rect 16686 4326 16698 4378
rect 16750 4326 16762 4378
rect 16814 4326 16826 4378
rect 16878 4326 16890 4378
rect 16942 4326 24476 4378
rect 24528 4326 24540 4378
rect 24592 4326 24604 4378
rect 24656 4326 24668 4378
rect 24720 4326 24732 4378
rect 24784 4326 32318 4378
rect 32370 4326 32382 4378
rect 32434 4326 32446 4378
rect 32498 4326 32510 4378
rect 32562 4326 32574 4378
rect 32626 4326 32632 4378
rect 1104 4304 32632 4326
rect 1104 3834 32476 3856
rect 1104 3782 4871 3834
rect 4923 3782 4935 3834
rect 4987 3782 4999 3834
rect 5051 3782 5063 3834
rect 5115 3782 5127 3834
rect 5179 3782 12713 3834
rect 12765 3782 12777 3834
rect 12829 3782 12841 3834
rect 12893 3782 12905 3834
rect 12957 3782 12969 3834
rect 13021 3782 20555 3834
rect 20607 3782 20619 3834
rect 20671 3782 20683 3834
rect 20735 3782 20747 3834
rect 20799 3782 20811 3834
rect 20863 3782 28397 3834
rect 28449 3782 28461 3834
rect 28513 3782 28525 3834
rect 28577 3782 28589 3834
rect 28641 3782 28653 3834
rect 28705 3782 32476 3834
rect 1104 3760 32476 3782
rect 1104 3290 32632 3312
rect 1104 3238 8792 3290
rect 8844 3238 8856 3290
rect 8908 3238 8920 3290
rect 8972 3238 8984 3290
rect 9036 3238 9048 3290
rect 9100 3238 16634 3290
rect 16686 3238 16698 3290
rect 16750 3238 16762 3290
rect 16814 3238 16826 3290
rect 16878 3238 16890 3290
rect 16942 3238 24476 3290
rect 24528 3238 24540 3290
rect 24592 3238 24604 3290
rect 24656 3238 24668 3290
rect 24720 3238 24732 3290
rect 24784 3238 32318 3290
rect 32370 3238 32382 3290
rect 32434 3238 32446 3290
rect 32498 3238 32510 3290
rect 32562 3238 32574 3290
rect 32626 3238 32632 3290
rect 1104 3216 32632 3238
rect 1104 2746 32476 2768
rect 1104 2694 4871 2746
rect 4923 2694 4935 2746
rect 4987 2694 4999 2746
rect 5051 2694 5063 2746
rect 5115 2694 5127 2746
rect 5179 2694 12713 2746
rect 12765 2694 12777 2746
rect 12829 2694 12841 2746
rect 12893 2694 12905 2746
rect 12957 2694 12969 2746
rect 13021 2694 20555 2746
rect 20607 2694 20619 2746
rect 20671 2694 20683 2746
rect 20735 2694 20747 2746
rect 20799 2694 20811 2746
rect 20863 2694 28397 2746
rect 28449 2694 28461 2746
rect 28513 2694 28525 2746
rect 28577 2694 28589 2746
rect 28641 2694 28653 2746
rect 28705 2694 32476 2746
rect 1104 2672 32476 2694
rect 1104 2202 32632 2224
rect 1104 2150 8792 2202
rect 8844 2150 8856 2202
rect 8908 2150 8920 2202
rect 8972 2150 8984 2202
rect 9036 2150 9048 2202
rect 9100 2150 16634 2202
rect 16686 2150 16698 2202
rect 16750 2150 16762 2202
rect 16814 2150 16826 2202
rect 16878 2150 16890 2202
rect 16942 2150 24476 2202
rect 24528 2150 24540 2202
rect 24592 2150 24604 2202
rect 24656 2150 24668 2202
rect 24720 2150 24732 2202
rect 24784 2150 32318 2202
rect 32370 2150 32382 2202
rect 32434 2150 32446 2202
rect 32498 2150 32510 2202
rect 32562 2150 32574 2202
rect 32626 2150 32632 2202
rect 1104 2128 32632 2150
rect 1104 1658 32476 1680
rect 1104 1606 4871 1658
rect 4923 1606 4935 1658
rect 4987 1606 4999 1658
rect 5051 1606 5063 1658
rect 5115 1606 5127 1658
rect 5179 1606 12713 1658
rect 12765 1606 12777 1658
rect 12829 1606 12841 1658
rect 12893 1606 12905 1658
rect 12957 1606 12969 1658
rect 13021 1606 20555 1658
rect 20607 1606 20619 1658
rect 20671 1606 20683 1658
rect 20735 1606 20747 1658
rect 20799 1606 20811 1658
rect 20863 1606 28397 1658
rect 28449 1606 28461 1658
rect 28513 1606 28525 1658
rect 28577 1606 28589 1658
rect 28641 1606 28653 1658
rect 28705 1606 32476 1658
rect 1104 1584 32476 1606
rect 1104 1114 32632 1136
rect 1104 1062 8792 1114
rect 8844 1062 8856 1114
rect 8908 1062 8920 1114
rect 8972 1062 8984 1114
rect 9036 1062 9048 1114
rect 9100 1062 16634 1114
rect 16686 1062 16698 1114
rect 16750 1062 16762 1114
rect 16814 1062 16826 1114
rect 16878 1062 16890 1114
rect 16942 1062 24476 1114
rect 24528 1062 24540 1114
rect 24592 1062 24604 1114
rect 24656 1062 24668 1114
rect 24720 1062 24732 1114
rect 24784 1062 32318 1114
rect 32370 1062 32382 1114
rect 32434 1062 32446 1114
rect 32498 1062 32510 1114
rect 32562 1062 32574 1114
rect 32626 1062 32632 1114
rect 1104 1040 32632 1062
<< via1 >>
rect 21552 21216 21612 21274
rect 33614 21208 33696 21280
rect 21732 21088 21784 21140
rect 24032 21088 24084 21140
rect 18420 21020 18472 21072
rect 19892 21020 19944 21072
rect 24124 21020 24176 21072
rect 18236 20952 18288 21004
rect 23112 20952 23164 21004
rect 19248 20884 19300 20936
rect 21088 20884 21140 20936
rect 19800 20816 19852 20868
rect 22468 20816 22520 20868
rect 28448 20816 28500 20868
rect 18052 20748 18104 20800
rect 22192 20748 22244 20800
rect 8792 20646 8844 20698
rect 8856 20646 8908 20698
rect 8920 20646 8972 20698
rect 8984 20646 9036 20698
rect 9048 20646 9100 20698
rect 16634 20646 16686 20698
rect 16698 20646 16750 20698
rect 16762 20646 16814 20698
rect 16826 20646 16878 20698
rect 16890 20646 16942 20698
rect 24476 20646 24528 20698
rect 24540 20646 24592 20698
rect 24604 20646 24656 20698
rect 24668 20646 24720 20698
rect 24732 20646 24784 20698
rect 32318 20646 32370 20698
rect 32382 20646 32434 20698
rect 32446 20646 32498 20698
rect 32510 20646 32562 20698
rect 32574 20646 32626 20698
rect 13820 20544 13872 20596
rect 2136 20451 2188 20460
rect 2136 20417 2145 20451
rect 2145 20417 2179 20451
rect 2179 20417 2188 20451
rect 2136 20408 2188 20417
rect 2780 20451 2832 20460
rect 2780 20417 2789 20451
rect 2789 20417 2823 20451
rect 2823 20417 2832 20451
rect 2780 20408 2832 20417
rect 3424 20451 3476 20460
rect 3424 20417 3433 20451
rect 3433 20417 3467 20451
rect 3467 20417 3476 20451
rect 3424 20408 3476 20417
rect 4528 20451 4580 20460
rect 4528 20417 4537 20451
rect 4537 20417 4571 20451
rect 4571 20417 4580 20451
rect 4528 20408 4580 20417
rect 5172 20451 5224 20460
rect 5172 20417 5181 20451
rect 5181 20417 5215 20451
rect 5215 20417 5224 20451
rect 5172 20408 5224 20417
rect 6000 20451 6052 20460
rect 6000 20417 6009 20451
rect 6009 20417 6043 20451
rect 6043 20417 6052 20451
rect 6000 20408 6052 20417
rect 7564 20451 7616 20460
rect 7564 20417 7573 20451
rect 7573 20417 7607 20451
rect 7607 20417 7616 20451
rect 7564 20408 7616 20417
rect 10232 20451 10284 20460
rect 10232 20417 10241 20451
rect 10241 20417 10275 20451
rect 10275 20417 10284 20451
rect 10232 20408 10284 20417
rect 12532 20476 12584 20528
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12440 20408 12492 20417
rect 14004 20476 14056 20528
rect 22284 20544 22336 20596
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 18236 20408 18288 20417
rect 19524 20408 19576 20460
rect 20168 20408 20220 20460
rect 20260 20451 20312 20460
rect 20260 20417 20269 20451
rect 20269 20417 20303 20451
rect 20303 20417 20312 20451
rect 20260 20408 20312 20417
rect 20352 20408 20404 20460
rect 22652 20476 22704 20528
rect 18144 20340 18196 20392
rect 21180 20340 21232 20392
rect 21916 20340 21968 20392
rect 22376 20451 22428 20460
rect 22376 20417 22385 20451
rect 22385 20417 22419 20451
rect 22419 20417 22428 20451
rect 22376 20408 22428 20417
rect 22744 20340 22796 20392
rect 12808 20272 12860 20324
rect 19892 20272 19944 20324
rect 20168 20272 20220 20324
rect 20996 20272 21048 20324
rect 23756 20544 23808 20596
rect 23848 20587 23900 20596
rect 23848 20553 23857 20587
rect 23857 20553 23891 20587
rect 23891 20553 23900 20587
rect 23848 20544 23900 20553
rect 24308 20544 24360 20596
rect 28448 20587 28500 20596
rect 28448 20553 28457 20587
rect 28457 20553 28491 20587
rect 28491 20553 28500 20587
rect 28448 20544 28500 20553
rect 23664 20476 23716 20528
rect 23572 20408 23624 20460
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 24216 20408 24268 20460
rect 25872 20408 25924 20460
rect 27344 20451 27396 20460
rect 27344 20417 27353 20451
rect 27353 20417 27387 20451
rect 27387 20417 27396 20451
rect 27344 20408 27396 20417
rect 27436 20408 27488 20460
rect 28632 20451 28684 20460
rect 28632 20417 28641 20451
rect 28641 20417 28675 20451
rect 28675 20417 28684 20451
rect 28632 20408 28684 20417
rect 29920 20451 29972 20460
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 30288 20408 30340 20460
rect 23388 20383 23440 20392
rect 23388 20349 23397 20383
rect 23397 20349 23431 20383
rect 23431 20349 23440 20383
rect 23388 20340 23440 20349
rect 24492 20340 24544 20392
rect 23480 20272 23532 20324
rect 11428 20204 11480 20256
rect 18880 20247 18932 20256
rect 18880 20213 18889 20247
rect 18889 20213 18923 20247
rect 18923 20213 18932 20247
rect 18880 20204 18932 20213
rect 20260 20204 20312 20256
rect 24860 20204 24912 20256
rect 25136 20247 25188 20256
rect 25136 20213 25145 20247
rect 25145 20213 25179 20247
rect 25179 20213 25188 20247
rect 25136 20204 25188 20213
rect 27160 20247 27212 20256
rect 27160 20213 27169 20247
rect 27169 20213 27203 20247
rect 27203 20213 27212 20247
rect 27160 20204 27212 20213
rect 27804 20247 27856 20256
rect 27804 20213 27813 20247
rect 27813 20213 27847 20247
rect 27847 20213 27856 20247
rect 27804 20204 27856 20213
rect 30380 20247 30432 20256
rect 30380 20213 30389 20247
rect 30389 20213 30423 20247
rect 30423 20213 30432 20247
rect 30380 20204 30432 20213
rect 4871 20102 4923 20154
rect 4935 20102 4987 20154
rect 4999 20102 5051 20154
rect 5063 20102 5115 20154
rect 5127 20102 5179 20154
rect 12713 20102 12765 20154
rect 12777 20102 12829 20154
rect 12841 20102 12893 20154
rect 12905 20102 12957 20154
rect 12969 20102 13021 20154
rect 20555 20102 20607 20154
rect 20619 20102 20671 20154
rect 20683 20102 20735 20154
rect 20747 20102 20799 20154
rect 20811 20102 20863 20154
rect 28397 20102 28449 20154
rect 28461 20102 28513 20154
rect 28525 20102 28577 20154
rect 28589 20102 28641 20154
rect 28653 20102 28705 20154
rect 1584 20043 1636 20052
rect 1584 20009 1593 20043
rect 1593 20009 1627 20043
rect 1627 20009 1636 20043
rect 1584 20000 1636 20009
rect 6736 20043 6788 20052
rect 6736 20009 6745 20043
rect 6745 20009 6779 20043
rect 6779 20009 6788 20043
rect 6736 20000 6788 20009
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 8208 20043 8260 20052
rect 8208 20009 8217 20043
rect 8217 20009 8251 20043
rect 8251 20009 8260 20043
rect 8208 20000 8260 20009
rect 9680 20000 9732 20052
rect 10140 20043 10192 20052
rect 10140 20009 10149 20043
rect 10149 20009 10183 20043
rect 10183 20009 10192 20043
rect 10140 20000 10192 20009
rect 11060 20000 11112 20052
rect 12624 20000 12676 20052
rect 17868 20000 17920 20052
rect 18420 20000 18472 20052
rect 18880 20000 18932 20052
rect 7564 19932 7616 19984
rect 15752 19932 15804 19984
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 12532 19864 12584 19916
rect 20812 19932 20864 19984
rect 21088 19932 21140 19984
rect 17224 19864 17276 19916
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 18052 19796 18104 19848
rect 19248 19796 19300 19848
rect 20352 19796 20404 19848
rect 20444 19796 20496 19848
rect 21548 19839 21600 19848
rect 21548 19805 21557 19839
rect 21557 19805 21591 19839
rect 21591 19805 21600 19839
rect 21548 19796 21600 19805
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 19524 19728 19576 19780
rect 18052 19660 18104 19712
rect 19800 19771 19852 19780
rect 19800 19737 19809 19771
rect 19809 19737 19843 19771
rect 19843 19737 19852 19771
rect 19800 19728 19852 19737
rect 19984 19728 20036 19780
rect 22284 19907 22336 19916
rect 22284 19873 22293 19907
rect 22293 19873 22327 19907
rect 22327 19873 22336 19907
rect 22284 19864 22336 19873
rect 23388 20000 23440 20052
rect 22836 19932 22888 19984
rect 22836 19796 22888 19848
rect 23480 19932 23532 19984
rect 23940 19932 23992 19984
rect 27804 19932 27856 19984
rect 24400 19864 24452 19916
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 28816 19796 28868 19848
rect 21640 19660 21692 19712
rect 23572 19728 23624 19780
rect 23296 19660 23348 19712
rect 25412 19703 25464 19712
rect 25412 19669 25421 19703
rect 25421 19669 25455 19703
rect 25455 19669 25464 19703
rect 25412 19660 25464 19669
rect 8792 19558 8844 19610
rect 8856 19558 8908 19610
rect 8920 19558 8972 19610
rect 8984 19558 9036 19610
rect 9048 19558 9100 19610
rect 16634 19558 16686 19610
rect 16698 19558 16750 19610
rect 16762 19558 16814 19610
rect 16826 19558 16878 19610
rect 16890 19558 16942 19610
rect 24476 19558 24528 19610
rect 24540 19558 24592 19610
rect 24604 19558 24656 19610
rect 24668 19558 24720 19610
rect 24732 19558 24784 19610
rect 32318 19558 32370 19610
rect 32382 19558 32434 19610
rect 32446 19558 32498 19610
rect 32510 19558 32562 19610
rect 32574 19558 32626 19610
rect 11428 19456 11480 19508
rect 17224 19456 17276 19508
rect 18052 19456 18104 19508
rect 19892 19456 19944 19508
rect 19800 19388 19852 19440
rect 22008 19456 22060 19508
rect 22100 19456 22152 19508
rect 22744 19456 22796 19508
rect 23020 19456 23072 19508
rect 27160 19456 27212 19508
rect 9128 19252 9180 19304
rect 11888 19295 11940 19304
rect 11888 19261 11897 19295
rect 11897 19261 11931 19295
rect 11931 19261 11940 19295
rect 11888 19252 11940 19261
rect 20904 19320 20956 19372
rect 19984 19252 20036 19304
rect 20628 19252 20680 19304
rect 10232 19184 10284 19236
rect 17224 19184 17276 19236
rect 17500 19227 17552 19236
rect 17500 19193 17509 19227
rect 17509 19193 17543 19227
rect 17543 19193 17552 19227
rect 17500 19184 17552 19193
rect 21456 19252 21508 19304
rect 21640 19252 21692 19304
rect 22468 19320 22520 19372
rect 22744 19252 22796 19304
rect 23296 19388 23348 19440
rect 23664 19388 23716 19440
rect 23388 19320 23440 19372
rect 23296 19252 23348 19304
rect 24216 19320 24268 19372
rect 22192 19184 22244 19236
rect 23756 19252 23808 19304
rect 24860 19320 24912 19372
rect 24216 19184 24268 19236
rect 21456 19116 21508 19168
rect 22284 19116 22336 19168
rect 23020 19116 23072 19168
rect 4871 19014 4923 19066
rect 4935 19014 4987 19066
rect 4999 19014 5051 19066
rect 5063 19014 5115 19066
rect 5127 19014 5179 19066
rect 12713 19014 12765 19066
rect 12777 19014 12829 19066
rect 12841 19014 12893 19066
rect 12905 19014 12957 19066
rect 12969 19014 13021 19066
rect 20555 19014 20607 19066
rect 20619 19014 20671 19066
rect 20683 19014 20735 19066
rect 20747 19014 20799 19066
rect 20811 19014 20863 19066
rect 28397 19014 28449 19066
rect 28461 19014 28513 19066
rect 28525 19014 28577 19066
rect 28589 19014 28641 19066
rect 28653 19014 28705 19066
rect 15568 18955 15620 18964
rect 15568 18921 15577 18955
rect 15577 18921 15611 18955
rect 15611 18921 15620 18955
rect 15568 18912 15620 18921
rect 22744 18955 22796 18964
rect 22744 18921 22753 18955
rect 22753 18921 22787 18955
rect 22787 18921 22796 18955
rect 22744 18912 22796 18921
rect 17224 18844 17276 18896
rect 17960 18819 18012 18828
rect 17960 18785 17969 18819
rect 17969 18785 18003 18819
rect 18003 18785 18012 18819
rect 17960 18776 18012 18785
rect 23112 18776 23164 18828
rect 17040 18751 17092 18760
rect 17040 18717 17049 18751
rect 17049 18717 17083 18751
rect 17083 18717 17092 18751
rect 17040 18708 17092 18717
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 22100 18751 22152 18760
rect 22100 18717 22109 18751
rect 22109 18717 22143 18751
rect 22143 18717 22152 18751
rect 22100 18708 22152 18717
rect 22284 18751 22336 18760
rect 22284 18717 22293 18751
rect 22293 18717 22327 18751
rect 22327 18717 22336 18751
rect 22284 18708 22336 18717
rect 22928 18751 22980 18760
rect 22928 18717 22937 18751
rect 22937 18717 22971 18751
rect 22971 18717 22980 18751
rect 22928 18708 22980 18717
rect 23480 18708 23532 18760
rect 23756 18708 23808 18760
rect 21916 18640 21968 18692
rect 24216 18640 24268 18692
rect 23480 18572 23532 18624
rect 8792 18470 8844 18522
rect 8856 18470 8908 18522
rect 8920 18470 8972 18522
rect 8984 18470 9036 18522
rect 9048 18470 9100 18522
rect 16634 18470 16686 18522
rect 16698 18470 16750 18522
rect 16762 18470 16814 18522
rect 16826 18470 16878 18522
rect 16890 18470 16942 18522
rect 24476 18470 24528 18522
rect 24540 18470 24592 18522
rect 24604 18470 24656 18522
rect 24668 18470 24720 18522
rect 24732 18470 24784 18522
rect 32318 18470 32370 18522
rect 32382 18470 32434 18522
rect 32446 18470 32498 18522
rect 32510 18470 32562 18522
rect 32574 18470 32626 18522
rect 23572 18411 23624 18420
rect 23572 18377 23581 18411
rect 23581 18377 23615 18411
rect 23615 18377 23624 18411
rect 23572 18368 23624 18377
rect 17040 18300 17092 18352
rect 25320 18300 25372 18352
rect 24032 18232 24084 18284
rect 4871 17926 4923 17978
rect 4935 17926 4987 17978
rect 4999 17926 5051 17978
rect 5063 17926 5115 17978
rect 5127 17926 5179 17978
rect 12713 17926 12765 17978
rect 12777 17926 12829 17978
rect 12841 17926 12893 17978
rect 12905 17926 12957 17978
rect 12969 17926 13021 17978
rect 20555 17926 20607 17978
rect 20619 17926 20671 17978
rect 20683 17926 20735 17978
rect 20747 17926 20799 17978
rect 20811 17926 20863 17978
rect 28397 17926 28449 17978
rect 28461 17926 28513 17978
rect 28525 17926 28577 17978
rect 28589 17926 28641 17978
rect 28653 17926 28705 17978
rect 22652 17824 22704 17876
rect 23480 17867 23532 17876
rect 23480 17833 23489 17867
rect 23489 17833 23523 17867
rect 23523 17833 23532 17867
rect 23480 17824 23532 17833
rect 23572 17688 23624 17740
rect 23940 17688 23992 17740
rect 23848 17620 23900 17672
rect 8792 17382 8844 17434
rect 8856 17382 8908 17434
rect 8920 17382 8972 17434
rect 8984 17382 9036 17434
rect 9048 17382 9100 17434
rect 16634 17382 16686 17434
rect 16698 17382 16750 17434
rect 16762 17382 16814 17434
rect 16826 17382 16878 17434
rect 16890 17382 16942 17434
rect 24476 17382 24528 17434
rect 24540 17382 24592 17434
rect 24604 17382 24656 17434
rect 24668 17382 24720 17434
rect 24732 17382 24784 17434
rect 32318 17382 32370 17434
rect 32382 17382 32434 17434
rect 32446 17382 32498 17434
rect 32510 17382 32562 17434
rect 32574 17382 32626 17434
rect 23664 17280 23716 17332
rect 19524 17144 19576 17196
rect 22376 17187 22428 17196
rect 22376 17153 22385 17187
rect 22385 17153 22419 17187
rect 22419 17153 22428 17187
rect 22376 17144 22428 17153
rect 22652 17144 22704 17196
rect 25136 17212 25188 17264
rect 23940 17144 23992 17196
rect 24124 17144 24176 17196
rect 23112 17119 23164 17128
rect 23112 17085 23121 17119
rect 23121 17085 23155 17119
rect 23155 17085 23164 17119
rect 23112 17076 23164 17085
rect 4871 16838 4923 16890
rect 4935 16838 4987 16890
rect 4999 16838 5051 16890
rect 5063 16838 5115 16890
rect 5127 16838 5179 16890
rect 12713 16838 12765 16890
rect 12777 16838 12829 16890
rect 12841 16838 12893 16890
rect 12905 16838 12957 16890
rect 12969 16838 13021 16890
rect 20555 16838 20607 16890
rect 20619 16838 20671 16890
rect 20683 16838 20735 16890
rect 20747 16838 20799 16890
rect 20811 16838 20863 16890
rect 28397 16838 28449 16890
rect 28461 16838 28513 16890
rect 28525 16838 28577 16890
rect 28589 16838 28641 16890
rect 28653 16838 28705 16890
rect 22376 16736 22428 16788
rect 24308 16600 24360 16652
rect 23848 16532 23900 16584
rect 23572 16507 23624 16516
rect 23572 16473 23581 16507
rect 23581 16473 23615 16507
rect 23615 16473 23624 16507
rect 23572 16464 23624 16473
rect 24124 16464 24176 16516
rect 24400 16464 24452 16516
rect 24032 16396 24084 16448
rect 8792 16294 8844 16346
rect 8856 16294 8908 16346
rect 8920 16294 8972 16346
rect 8984 16294 9036 16346
rect 9048 16294 9100 16346
rect 16634 16294 16686 16346
rect 16698 16294 16750 16346
rect 16762 16294 16814 16346
rect 16826 16294 16878 16346
rect 16890 16294 16942 16346
rect 24476 16294 24528 16346
rect 24540 16294 24592 16346
rect 24604 16294 24656 16346
rect 24668 16294 24720 16346
rect 24732 16294 24784 16346
rect 32318 16294 32370 16346
rect 32382 16294 32434 16346
rect 32446 16294 32498 16346
rect 32510 16294 32562 16346
rect 32574 16294 32626 16346
rect 17868 16192 17920 16244
rect 20996 16056 21048 16108
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 18052 15920 18104 15972
rect 4871 15750 4923 15802
rect 4935 15750 4987 15802
rect 4999 15750 5051 15802
rect 5063 15750 5115 15802
rect 5127 15750 5179 15802
rect 12713 15750 12765 15802
rect 12777 15750 12829 15802
rect 12841 15750 12893 15802
rect 12905 15750 12957 15802
rect 12969 15750 13021 15802
rect 20555 15750 20607 15802
rect 20619 15750 20671 15802
rect 20683 15750 20735 15802
rect 20747 15750 20799 15802
rect 20811 15750 20863 15802
rect 28397 15750 28449 15802
rect 28461 15750 28513 15802
rect 28525 15750 28577 15802
rect 28589 15750 28641 15802
rect 28653 15750 28705 15802
rect 8792 15206 8844 15258
rect 8856 15206 8908 15258
rect 8920 15206 8972 15258
rect 8984 15206 9036 15258
rect 9048 15206 9100 15258
rect 16634 15206 16686 15258
rect 16698 15206 16750 15258
rect 16762 15206 16814 15258
rect 16826 15206 16878 15258
rect 16890 15206 16942 15258
rect 24476 15206 24528 15258
rect 24540 15206 24592 15258
rect 24604 15206 24656 15258
rect 24668 15206 24720 15258
rect 24732 15206 24784 15258
rect 32318 15206 32370 15258
rect 32382 15206 32434 15258
rect 32446 15206 32498 15258
rect 32510 15206 32562 15258
rect 32574 15206 32626 15258
rect 21548 15104 21600 15156
rect 25320 15104 25372 15156
rect 23940 15036 23992 15088
rect 24124 14968 24176 15020
rect 24400 14968 24452 15020
rect 25136 14968 25188 15020
rect 23664 14900 23716 14952
rect 4871 14662 4923 14714
rect 4935 14662 4987 14714
rect 4999 14662 5051 14714
rect 5063 14662 5115 14714
rect 5127 14662 5179 14714
rect 12713 14662 12765 14714
rect 12777 14662 12829 14714
rect 12841 14662 12893 14714
rect 12905 14662 12957 14714
rect 12969 14662 13021 14714
rect 20555 14662 20607 14714
rect 20619 14662 20671 14714
rect 20683 14662 20735 14714
rect 20747 14662 20799 14714
rect 20811 14662 20863 14714
rect 28397 14662 28449 14714
rect 28461 14662 28513 14714
rect 28525 14662 28577 14714
rect 28589 14662 28641 14714
rect 28653 14662 28705 14714
rect 20444 14560 20496 14612
rect 19800 14424 19852 14476
rect 20168 14467 20220 14476
rect 20168 14433 20177 14467
rect 20177 14433 20211 14467
rect 20211 14433 20220 14467
rect 20168 14424 20220 14433
rect 25504 14356 25556 14408
rect 8792 14118 8844 14170
rect 8856 14118 8908 14170
rect 8920 14118 8972 14170
rect 8984 14118 9036 14170
rect 9048 14118 9100 14170
rect 16634 14118 16686 14170
rect 16698 14118 16750 14170
rect 16762 14118 16814 14170
rect 16826 14118 16878 14170
rect 16890 14118 16942 14170
rect 24476 14118 24528 14170
rect 24540 14118 24592 14170
rect 24604 14118 24656 14170
rect 24668 14118 24720 14170
rect 24732 14118 24784 14170
rect 32318 14118 32370 14170
rect 32382 14118 32434 14170
rect 32446 14118 32498 14170
rect 32510 14118 32562 14170
rect 32574 14118 32626 14170
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 20168 13948 20220 14000
rect 25412 13948 25464 14000
rect 30380 13948 30432 14000
rect 4871 13574 4923 13626
rect 4935 13574 4987 13626
rect 4999 13574 5051 13626
rect 5063 13574 5115 13626
rect 5127 13574 5179 13626
rect 12713 13574 12765 13626
rect 12777 13574 12829 13626
rect 12841 13574 12893 13626
rect 12905 13574 12957 13626
rect 12969 13574 13021 13626
rect 20555 13574 20607 13626
rect 20619 13574 20671 13626
rect 20683 13574 20735 13626
rect 20747 13574 20799 13626
rect 20811 13574 20863 13626
rect 28397 13574 28449 13626
rect 28461 13574 28513 13626
rect 28525 13574 28577 13626
rect 28589 13574 28641 13626
rect 28653 13574 28705 13626
rect 8792 13030 8844 13082
rect 8856 13030 8908 13082
rect 8920 13030 8972 13082
rect 8984 13030 9036 13082
rect 9048 13030 9100 13082
rect 16634 13030 16686 13082
rect 16698 13030 16750 13082
rect 16762 13030 16814 13082
rect 16826 13030 16878 13082
rect 16890 13030 16942 13082
rect 24476 13030 24528 13082
rect 24540 13030 24592 13082
rect 24604 13030 24656 13082
rect 24668 13030 24720 13082
rect 24732 13030 24784 13082
rect 32318 13030 32370 13082
rect 32382 13030 32434 13082
rect 32446 13030 32498 13082
rect 32510 13030 32562 13082
rect 32574 13030 32626 13082
rect 23756 12792 23808 12844
rect 12440 12588 12492 12640
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 4871 12486 4923 12538
rect 4935 12486 4987 12538
rect 4999 12486 5051 12538
rect 5063 12486 5115 12538
rect 5127 12486 5179 12538
rect 12713 12486 12765 12538
rect 12777 12486 12829 12538
rect 12841 12486 12893 12538
rect 12905 12486 12957 12538
rect 12969 12486 13021 12538
rect 20555 12486 20607 12538
rect 20619 12486 20671 12538
rect 20683 12486 20735 12538
rect 20747 12486 20799 12538
rect 20811 12486 20863 12538
rect 28397 12486 28449 12538
rect 28461 12486 28513 12538
rect 28525 12486 28577 12538
rect 28589 12486 28641 12538
rect 28653 12486 28705 12538
rect 20996 12384 21048 12436
rect 21640 12384 21692 12436
rect 24032 12248 24084 12300
rect 20168 12112 20220 12164
rect 8792 11942 8844 11994
rect 8856 11942 8908 11994
rect 8920 11942 8972 11994
rect 8984 11942 9036 11994
rect 9048 11942 9100 11994
rect 16634 11942 16686 11994
rect 16698 11942 16750 11994
rect 16762 11942 16814 11994
rect 16826 11942 16878 11994
rect 16890 11942 16942 11994
rect 24476 11942 24528 11994
rect 24540 11942 24592 11994
rect 24604 11942 24656 11994
rect 24668 11942 24720 11994
rect 24732 11942 24784 11994
rect 32318 11942 32370 11994
rect 32382 11942 32434 11994
rect 32446 11942 32498 11994
rect 32510 11942 32562 11994
rect 32574 11942 32626 11994
rect 4871 11398 4923 11450
rect 4935 11398 4987 11450
rect 4999 11398 5051 11450
rect 5063 11398 5115 11450
rect 5127 11398 5179 11450
rect 12713 11398 12765 11450
rect 12777 11398 12829 11450
rect 12841 11398 12893 11450
rect 12905 11398 12957 11450
rect 12969 11398 13021 11450
rect 20555 11398 20607 11450
rect 20619 11398 20671 11450
rect 20683 11398 20735 11450
rect 20747 11398 20799 11450
rect 20811 11398 20863 11450
rect 28397 11398 28449 11450
rect 28461 11398 28513 11450
rect 28525 11398 28577 11450
rect 28589 11398 28641 11450
rect 28653 11398 28705 11450
rect 8792 10854 8844 10906
rect 8856 10854 8908 10906
rect 8920 10854 8972 10906
rect 8984 10854 9036 10906
rect 9048 10854 9100 10906
rect 16634 10854 16686 10906
rect 16698 10854 16750 10906
rect 16762 10854 16814 10906
rect 16826 10854 16878 10906
rect 16890 10854 16942 10906
rect 24476 10854 24528 10906
rect 24540 10854 24592 10906
rect 24604 10854 24656 10906
rect 24668 10854 24720 10906
rect 24732 10854 24784 10906
rect 32318 10854 32370 10906
rect 32382 10854 32434 10906
rect 32446 10854 32498 10906
rect 32510 10854 32562 10906
rect 32574 10854 32626 10906
rect 4871 10310 4923 10362
rect 4935 10310 4987 10362
rect 4999 10310 5051 10362
rect 5063 10310 5115 10362
rect 5127 10310 5179 10362
rect 12713 10310 12765 10362
rect 12777 10310 12829 10362
rect 12841 10310 12893 10362
rect 12905 10310 12957 10362
rect 12969 10310 13021 10362
rect 20555 10310 20607 10362
rect 20619 10310 20671 10362
rect 20683 10310 20735 10362
rect 20747 10310 20799 10362
rect 20811 10310 20863 10362
rect 28397 10310 28449 10362
rect 28461 10310 28513 10362
rect 28525 10310 28577 10362
rect 28589 10310 28641 10362
rect 28653 10310 28705 10362
rect 8792 9766 8844 9818
rect 8856 9766 8908 9818
rect 8920 9766 8972 9818
rect 8984 9766 9036 9818
rect 9048 9766 9100 9818
rect 16634 9766 16686 9818
rect 16698 9766 16750 9818
rect 16762 9766 16814 9818
rect 16826 9766 16878 9818
rect 16890 9766 16942 9818
rect 24476 9766 24528 9818
rect 24540 9766 24592 9818
rect 24604 9766 24656 9818
rect 24668 9766 24720 9818
rect 24732 9766 24784 9818
rect 32318 9766 32370 9818
rect 32382 9766 32434 9818
rect 32446 9766 32498 9818
rect 32510 9766 32562 9818
rect 32574 9766 32626 9818
rect 4871 9222 4923 9274
rect 4935 9222 4987 9274
rect 4999 9222 5051 9274
rect 5063 9222 5115 9274
rect 5127 9222 5179 9274
rect 12713 9222 12765 9274
rect 12777 9222 12829 9274
rect 12841 9222 12893 9274
rect 12905 9222 12957 9274
rect 12969 9222 13021 9274
rect 20555 9222 20607 9274
rect 20619 9222 20671 9274
rect 20683 9222 20735 9274
rect 20747 9222 20799 9274
rect 20811 9222 20863 9274
rect 28397 9222 28449 9274
rect 28461 9222 28513 9274
rect 28525 9222 28577 9274
rect 28589 9222 28641 9274
rect 28653 9222 28705 9274
rect 8792 8678 8844 8730
rect 8856 8678 8908 8730
rect 8920 8678 8972 8730
rect 8984 8678 9036 8730
rect 9048 8678 9100 8730
rect 16634 8678 16686 8730
rect 16698 8678 16750 8730
rect 16762 8678 16814 8730
rect 16826 8678 16878 8730
rect 16890 8678 16942 8730
rect 24476 8678 24528 8730
rect 24540 8678 24592 8730
rect 24604 8678 24656 8730
rect 24668 8678 24720 8730
rect 24732 8678 24784 8730
rect 32318 8678 32370 8730
rect 32382 8678 32434 8730
rect 32446 8678 32498 8730
rect 32510 8678 32562 8730
rect 32574 8678 32626 8730
rect 4871 8134 4923 8186
rect 4935 8134 4987 8186
rect 4999 8134 5051 8186
rect 5063 8134 5115 8186
rect 5127 8134 5179 8186
rect 12713 8134 12765 8186
rect 12777 8134 12829 8186
rect 12841 8134 12893 8186
rect 12905 8134 12957 8186
rect 12969 8134 13021 8186
rect 20555 8134 20607 8186
rect 20619 8134 20671 8186
rect 20683 8134 20735 8186
rect 20747 8134 20799 8186
rect 20811 8134 20863 8186
rect 28397 8134 28449 8186
rect 28461 8134 28513 8186
rect 28525 8134 28577 8186
rect 28589 8134 28641 8186
rect 28653 8134 28705 8186
rect 8792 7590 8844 7642
rect 8856 7590 8908 7642
rect 8920 7590 8972 7642
rect 8984 7590 9036 7642
rect 9048 7590 9100 7642
rect 16634 7590 16686 7642
rect 16698 7590 16750 7642
rect 16762 7590 16814 7642
rect 16826 7590 16878 7642
rect 16890 7590 16942 7642
rect 24476 7590 24528 7642
rect 24540 7590 24592 7642
rect 24604 7590 24656 7642
rect 24668 7590 24720 7642
rect 24732 7590 24784 7642
rect 32318 7590 32370 7642
rect 32382 7590 32434 7642
rect 32446 7590 32498 7642
rect 32510 7590 32562 7642
rect 32574 7590 32626 7642
rect 4871 7046 4923 7098
rect 4935 7046 4987 7098
rect 4999 7046 5051 7098
rect 5063 7046 5115 7098
rect 5127 7046 5179 7098
rect 12713 7046 12765 7098
rect 12777 7046 12829 7098
rect 12841 7046 12893 7098
rect 12905 7046 12957 7098
rect 12969 7046 13021 7098
rect 20555 7046 20607 7098
rect 20619 7046 20671 7098
rect 20683 7046 20735 7098
rect 20747 7046 20799 7098
rect 20811 7046 20863 7098
rect 28397 7046 28449 7098
rect 28461 7046 28513 7098
rect 28525 7046 28577 7098
rect 28589 7046 28641 7098
rect 28653 7046 28705 7098
rect 8792 6502 8844 6554
rect 8856 6502 8908 6554
rect 8920 6502 8972 6554
rect 8984 6502 9036 6554
rect 9048 6502 9100 6554
rect 16634 6502 16686 6554
rect 16698 6502 16750 6554
rect 16762 6502 16814 6554
rect 16826 6502 16878 6554
rect 16890 6502 16942 6554
rect 24476 6502 24528 6554
rect 24540 6502 24592 6554
rect 24604 6502 24656 6554
rect 24668 6502 24720 6554
rect 24732 6502 24784 6554
rect 32318 6502 32370 6554
rect 32382 6502 32434 6554
rect 32446 6502 32498 6554
rect 32510 6502 32562 6554
rect 32574 6502 32626 6554
rect 4871 5958 4923 6010
rect 4935 5958 4987 6010
rect 4999 5958 5051 6010
rect 5063 5958 5115 6010
rect 5127 5958 5179 6010
rect 12713 5958 12765 6010
rect 12777 5958 12829 6010
rect 12841 5958 12893 6010
rect 12905 5958 12957 6010
rect 12969 5958 13021 6010
rect 20555 5958 20607 6010
rect 20619 5958 20671 6010
rect 20683 5958 20735 6010
rect 20747 5958 20799 6010
rect 20811 5958 20863 6010
rect 28397 5958 28449 6010
rect 28461 5958 28513 6010
rect 28525 5958 28577 6010
rect 28589 5958 28641 6010
rect 28653 5958 28705 6010
rect 8792 5414 8844 5466
rect 8856 5414 8908 5466
rect 8920 5414 8972 5466
rect 8984 5414 9036 5466
rect 9048 5414 9100 5466
rect 16634 5414 16686 5466
rect 16698 5414 16750 5466
rect 16762 5414 16814 5466
rect 16826 5414 16878 5466
rect 16890 5414 16942 5466
rect 24476 5414 24528 5466
rect 24540 5414 24592 5466
rect 24604 5414 24656 5466
rect 24668 5414 24720 5466
rect 24732 5414 24784 5466
rect 32318 5414 32370 5466
rect 32382 5414 32434 5466
rect 32446 5414 32498 5466
rect 32510 5414 32562 5466
rect 32574 5414 32626 5466
rect 4871 4870 4923 4922
rect 4935 4870 4987 4922
rect 4999 4870 5051 4922
rect 5063 4870 5115 4922
rect 5127 4870 5179 4922
rect 12713 4870 12765 4922
rect 12777 4870 12829 4922
rect 12841 4870 12893 4922
rect 12905 4870 12957 4922
rect 12969 4870 13021 4922
rect 20555 4870 20607 4922
rect 20619 4870 20671 4922
rect 20683 4870 20735 4922
rect 20747 4870 20799 4922
rect 20811 4870 20863 4922
rect 28397 4870 28449 4922
rect 28461 4870 28513 4922
rect 28525 4870 28577 4922
rect 28589 4870 28641 4922
rect 28653 4870 28705 4922
rect 8792 4326 8844 4378
rect 8856 4326 8908 4378
rect 8920 4326 8972 4378
rect 8984 4326 9036 4378
rect 9048 4326 9100 4378
rect 16634 4326 16686 4378
rect 16698 4326 16750 4378
rect 16762 4326 16814 4378
rect 16826 4326 16878 4378
rect 16890 4326 16942 4378
rect 24476 4326 24528 4378
rect 24540 4326 24592 4378
rect 24604 4326 24656 4378
rect 24668 4326 24720 4378
rect 24732 4326 24784 4378
rect 32318 4326 32370 4378
rect 32382 4326 32434 4378
rect 32446 4326 32498 4378
rect 32510 4326 32562 4378
rect 32574 4326 32626 4378
rect 4871 3782 4923 3834
rect 4935 3782 4987 3834
rect 4999 3782 5051 3834
rect 5063 3782 5115 3834
rect 5127 3782 5179 3834
rect 12713 3782 12765 3834
rect 12777 3782 12829 3834
rect 12841 3782 12893 3834
rect 12905 3782 12957 3834
rect 12969 3782 13021 3834
rect 20555 3782 20607 3834
rect 20619 3782 20671 3834
rect 20683 3782 20735 3834
rect 20747 3782 20799 3834
rect 20811 3782 20863 3834
rect 28397 3782 28449 3834
rect 28461 3782 28513 3834
rect 28525 3782 28577 3834
rect 28589 3782 28641 3834
rect 28653 3782 28705 3834
rect 8792 3238 8844 3290
rect 8856 3238 8908 3290
rect 8920 3238 8972 3290
rect 8984 3238 9036 3290
rect 9048 3238 9100 3290
rect 16634 3238 16686 3290
rect 16698 3238 16750 3290
rect 16762 3238 16814 3290
rect 16826 3238 16878 3290
rect 16890 3238 16942 3290
rect 24476 3238 24528 3290
rect 24540 3238 24592 3290
rect 24604 3238 24656 3290
rect 24668 3238 24720 3290
rect 24732 3238 24784 3290
rect 32318 3238 32370 3290
rect 32382 3238 32434 3290
rect 32446 3238 32498 3290
rect 32510 3238 32562 3290
rect 32574 3238 32626 3290
rect 4871 2694 4923 2746
rect 4935 2694 4987 2746
rect 4999 2694 5051 2746
rect 5063 2694 5115 2746
rect 5127 2694 5179 2746
rect 12713 2694 12765 2746
rect 12777 2694 12829 2746
rect 12841 2694 12893 2746
rect 12905 2694 12957 2746
rect 12969 2694 13021 2746
rect 20555 2694 20607 2746
rect 20619 2694 20671 2746
rect 20683 2694 20735 2746
rect 20747 2694 20799 2746
rect 20811 2694 20863 2746
rect 28397 2694 28449 2746
rect 28461 2694 28513 2746
rect 28525 2694 28577 2746
rect 28589 2694 28641 2746
rect 28653 2694 28705 2746
rect 8792 2150 8844 2202
rect 8856 2150 8908 2202
rect 8920 2150 8972 2202
rect 8984 2150 9036 2202
rect 9048 2150 9100 2202
rect 16634 2150 16686 2202
rect 16698 2150 16750 2202
rect 16762 2150 16814 2202
rect 16826 2150 16878 2202
rect 16890 2150 16942 2202
rect 24476 2150 24528 2202
rect 24540 2150 24592 2202
rect 24604 2150 24656 2202
rect 24668 2150 24720 2202
rect 24732 2150 24784 2202
rect 32318 2150 32370 2202
rect 32382 2150 32434 2202
rect 32446 2150 32498 2202
rect 32510 2150 32562 2202
rect 32574 2150 32626 2202
rect 4871 1606 4923 1658
rect 4935 1606 4987 1658
rect 4999 1606 5051 1658
rect 5063 1606 5115 1658
rect 5127 1606 5179 1658
rect 12713 1606 12765 1658
rect 12777 1606 12829 1658
rect 12841 1606 12893 1658
rect 12905 1606 12957 1658
rect 12969 1606 13021 1658
rect 20555 1606 20607 1658
rect 20619 1606 20671 1658
rect 20683 1606 20735 1658
rect 20747 1606 20799 1658
rect 20811 1606 20863 1658
rect 28397 1606 28449 1658
rect 28461 1606 28513 1658
rect 28525 1606 28577 1658
rect 28589 1606 28641 1658
rect 28653 1606 28705 1658
rect 8792 1062 8844 1114
rect 8856 1062 8908 1114
rect 8920 1062 8972 1114
rect 8984 1062 9036 1114
rect 9048 1062 9100 1114
rect 16634 1062 16686 1114
rect 16698 1062 16750 1114
rect 16762 1062 16814 1114
rect 16826 1062 16878 1114
rect 16890 1062 16942 1114
rect 24476 1062 24528 1114
rect 24540 1062 24592 1114
rect 24604 1062 24656 1114
rect 24668 1062 24720 1114
rect 24732 1062 24784 1114
rect 32318 1062 32370 1114
rect 32382 1062 32434 1114
rect 32446 1062 32498 1114
rect 32510 1062 32562 1114
rect 32574 1062 32626 1114
<< metal2 >>
rect 9126 21448 9182 21457
rect 9126 21383 9182 21392
rect 9678 21448 9734 21457
rect 9678 21383 9734 21392
rect 11058 21448 11114 21457
rect 11058 21383 11114 21392
rect 11886 21448 11942 21457
rect 11886 21383 11942 21392
rect 12806 21448 12862 21457
rect 12806 21383 12862 21392
rect 14002 21448 14058 21457
rect 14002 21383 14058 21392
rect 15566 21448 15622 21457
rect 15566 21383 15622 21392
rect 15750 21448 15806 21457
rect 15750 21383 15806 21392
rect 17498 21448 17554 21457
rect 17498 21383 17554 21392
rect 19246 21448 19302 21457
rect 19246 21383 19302 21392
rect 19522 21448 19578 21457
rect 19522 21383 19578 21392
rect 21730 21448 21786 21457
rect 21730 21383 21786 21392
rect 22926 21448 22982 21457
rect 22926 21383 22982 21392
rect 23662 21448 23718 21457
rect 23662 21383 23718 21392
rect 24398 21448 24454 21457
rect 24398 21383 24454 21392
rect 25870 21448 25926 21457
rect 25870 21383 25926 21392
rect 27434 21448 27490 21457
rect 27434 21383 27490 21392
rect 28814 21448 28870 21457
rect 28814 21383 28870 21392
rect 30286 21448 30342 21457
rect 30286 21383 30342 21392
rect 5170 20904 5226 20913
rect 5170 20839 5226 20848
rect 2134 20496 2190 20505
rect 2134 20431 2136 20440
rect 2188 20431 2190 20440
rect 2778 20496 2834 20505
rect 2778 20431 2780 20440
rect 2136 20402 2188 20408
rect 2832 20431 2834 20440
rect 3422 20496 3478 20505
rect 3422 20431 3424 20440
rect 2780 20402 2832 20408
rect 3476 20431 3478 20440
rect 4526 20496 4582 20505
rect 5184 20466 5212 20839
rect 8792 20700 9100 20709
rect 8792 20698 8798 20700
rect 8854 20698 8878 20700
rect 8934 20698 8958 20700
rect 9014 20698 9038 20700
rect 9094 20698 9100 20700
rect 8854 20646 8856 20698
rect 9036 20646 9038 20698
rect 8792 20644 8798 20646
rect 8854 20644 8878 20646
rect 8934 20644 8958 20646
rect 9014 20644 9038 20646
rect 9094 20644 9100 20646
rect 8792 20635 9100 20644
rect 5998 20496 6054 20505
rect 4526 20431 4528 20440
rect 3424 20402 3476 20408
rect 4580 20431 4582 20440
rect 5172 20460 5224 20466
rect 4528 20402 4580 20408
rect 5998 20431 6000 20440
rect 5172 20402 5224 20408
rect 6052 20431 6054 20440
rect 7564 20460 7616 20466
rect 6000 20402 6052 20408
rect 7564 20402 7616 20408
rect 4871 20156 5179 20165
rect 4871 20154 4877 20156
rect 4933 20154 4957 20156
rect 5013 20154 5037 20156
rect 5093 20154 5117 20156
rect 5173 20154 5179 20156
rect 4933 20102 4935 20154
rect 5115 20102 5117 20154
rect 4871 20100 4877 20102
rect 4933 20100 4957 20102
rect 5013 20100 5037 20102
rect 5093 20100 5117 20102
rect 5173 20100 5179 20102
rect 1582 20088 1638 20097
rect 4871 20091 5179 20100
rect 1582 20023 1584 20032
rect 1636 20023 1638 20032
rect 6734 20088 6790 20097
rect 6734 20023 6736 20032
rect 1584 19994 1636 20000
rect 6788 20023 6790 20032
rect 7470 20088 7526 20097
rect 7470 20023 7472 20032
rect 6736 19994 6788 20000
rect 7524 20023 7526 20032
rect 7472 19994 7524 20000
rect 7576 19990 7604 20402
rect 8206 20088 8262 20097
rect 8206 20023 8208 20032
rect 8260 20023 8262 20032
rect 8208 19994 8260 20000
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 8792 19612 9100 19621
rect 8792 19610 8798 19612
rect 8854 19610 8878 19612
rect 8934 19610 8958 19612
rect 9014 19610 9038 19612
rect 9094 19610 9100 19612
rect 8854 19558 8856 19610
rect 9036 19558 9038 19610
rect 8792 19556 8798 19558
rect 8854 19556 8878 19558
rect 8934 19556 8958 19558
rect 9014 19556 9038 19558
rect 9094 19556 9100 19558
rect 8792 19547 9100 19556
rect 9140 19310 9168 21383
rect 9692 20058 9720 21383
rect 10232 20460 10284 20466
rect 10232 20402 10284 20408
rect 10138 20088 10194 20097
rect 9680 20052 9732 20058
rect 10138 20023 10140 20032
rect 9680 19994 9732 20000
rect 10192 20023 10194 20032
rect 10140 19994 10192 20000
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 10244 19242 10272 20402
rect 11072 20058 11100 21383
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11440 19854 11468 20198
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11440 19514 11468 19790
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11900 19310 11928 21383
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 10232 19236 10284 19242
rect 10232 19178 10284 19184
rect 4871 19068 5179 19077
rect 4871 19066 4877 19068
rect 4933 19066 4957 19068
rect 5013 19066 5037 19068
rect 5093 19066 5117 19068
rect 5173 19066 5179 19068
rect 4933 19014 4935 19066
rect 5115 19014 5117 19066
rect 4871 19012 4877 19014
rect 4933 19012 4957 19014
rect 5013 19012 5037 19014
rect 5093 19012 5117 19014
rect 5173 19012 5179 19014
rect 4871 19003 5179 19012
rect 8792 18524 9100 18533
rect 8792 18522 8798 18524
rect 8854 18522 8878 18524
rect 8934 18522 8958 18524
rect 9014 18522 9038 18524
rect 9094 18522 9100 18524
rect 8854 18470 8856 18522
rect 9036 18470 9038 18522
rect 8792 18468 8798 18470
rect 8854 18468 8878 18470
rect 8934 18468 8958 18470
rect 9014 18468 9038 18470
rect 9094 18468 9100 18470
rect 8792 18459 9100 18468
rect 4871 17980 5179 17989
rect 4871 17978 4877 17980
rect 4933 17978 4957 17980
rect 5013 17978 5037 17980
rect 5093 17978 5117 17980
rect 5173 17978 5179 17980
rect 4933 17926 4935 17978
rect 5115 17926 5117 17978
rect 4871 17924 4877 17926
rect 4933 17924 4957 17926
rect 5013 17924 5037 17926
rect 5093 17924 5117 17926
rect 5173 17924 5179 17926
rect 4871 17915 5179 17924
rect 8792 17436 9100 17445
rect 8792 17434 8798 17436
rect 8854 17434 8878 17436
rect 8934 17434 8958 17436
rect 9014 17434 9038 17436
rect 9094 17434 9100 17436
rect 8854 17382 8856 17434
rect 9036 17382 9038 17434
rect 8792 17380 8798 17382
rect 8854 17380 8878 17382
rect 8934 17380 8958 17382
rect 9014 17380 9038 17382
rect 9094 17380 9100 17382
rect 8792 17371 9100 17380
rect 4871 16892 5179 16901
rect 4871 16890 4877 16892
rect 4933 16890 4957 16892
rect 5013 16890 5037 16892
rect 5093 16890 5117 16892
rect 5173 16890 5179 16892
rect 4933 16838 4935 16890
rect 5115 16838 5117 16890
rect 4871 16836 4877 16838
rect 4933 16836 4957 16838
rect 5013 16836 5037 16838
rect 5093 16836 5117 16838
rect 5173 16836 5179 16838
rect 4871 16827 5179 16836
rect 8792 16348 9100 16357
rect 8792 16346 8798 16348
rect 8854 16346 8878 16348
rect 8934 16346 8958 16348
rect 9014 16346 9038 16348
rect 9094 16346 9100 16348
rect 8854 16294 8856 16346
rect 9036 16294 9038 16346
rect 8792 16292 8798 16294
rect 8854 16292 8878 16294
rect 8934 16292 8958 16294
rect 9014 16292 9038 16294
rect 9094 16292 9100 16294
rect 8792 16283 9100 16292
rect 4871 15804 5179 15813
rect 4871 15802 4877 15804
rect 4933 15802 4957 15804
rect 5013 15802 5037 15804
rect 5093 15802 5117 15804
rect 5173 15802 5179 15804
rect 4933 15750 4935 15802
rect 5115 15750 5117 15802
rect 4871 15748 4877 15750
rect 4933 15748 4957 15750
rect 5013 15748 5037 15750
rect 5093 15748 5117 15750
rect 5173 15748 5179 15750
rect 4871 15739 5179 15748
rect 8792 15260 9100 15269
rect 8792 15258 8798 15260
rect 8854 15258 8878 15260
rect 8934 15258 8958 15260
rect 9014 15258 9038 15260
rect 9094 15258 9100 15260
rect 8854 15206 8856 15258
rect 9036 15206 9038 15258
rect 8792 15204 8798 15206
rect 8854 15204 8878 15206
rect 8934 15204 8958 15206
rect 9014 15204 9038 15206
rect 9094 15204 9100 15206
rect 8792 15195 9100 15204
rect 4871 14716 5179 14725
rect 4871 14714 4877 14716
rect 4933 14714 4957 14716
rect 5013 14714 5037 14716
rect 5093 14714 5117 14716
rect 5173 14714 5179 14716
rect 4933 14662 4935 14714
rect 5115 14662 5117 14714
rect 4871 14660 4877 14662
rect 4933 14660 4957 14662
rect 5013 14660 5037 14662
rect 5093 14660 5117 14662
rect 5173 14660 5179 14662
rect 4871 14651 5179 14660
rect 8792 14172 9100 14181
rect 8792 14170 8798 14172
rect 8854 14170 8878 14172
rect 8934 14170 8958 14172
rect 9014 14170 9038 14172
rect 9094 14170 9100 14172
rect 8854 14118 8856 14170
rect 9036 14118 9038 14170
rect 8792 14116 8798 14118
rect 8854 14116 8878 14118
rect 8934 14116 8958 14118
rect 9014 14116 9038 14118
rect 9094 14116 9100 14118
rect 8792 14107 9100 14116
rect 4871 13628 5179 13637
rect 4871 13626 4877 13628
rect 4933 13626 4957 13628
rect 5013 13626 5037 13628
rect 5093 13626 5117 13628
rect 5173 13626 5179 13628
rect 4933 13574 4935 13626
rect 5115 13574 5117 13626
rect 4871 13572 4877 13574
rect 4933 13572 4957 13574
rect 5013 13572 5037 13574
rect 5093 13572 5117 13574
rect 5173 13572 5179 13574
rect 4871 13563 5179 13572
rect 8792 13084 9100 13093
rect 8792 13082 8798 13084
rect 8854 13082 8878 13084
rect 8934 13082 8958 13084
rect 9014 13082 9038 13084
rect 9094 13082 9100 13084
rect 8854 13030 8856 13082
rect 9036 13030 9038 13082
rect 8792 13028 8798 13030
rect 8854 13028 8878 13030
rect 8934 13028 8958 13030
rect 9014 13028 9038 13030
rect 9094 13028 9100 13030
rect 8792 13019 9100 13028
rect 12452 12646 12480 20402
rect 12544 19922 12572 20470
rect 12622 20360 12678 20369
rect 12820 20330 12848 21383
rect 13818 21312 13874 21321
rect 13818 21247 13874 21256
rect 13832 20602 13860 21247
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 14016 20534 14044 21383
rect 14004 20528 14056 20534
rect 14004 20470 14056 20476
rect 12622 20295 12678 20304
rect 12808 20324 12860 20330
rect 12636 20058 12664 20295
rect 12808 20266 12860 20272
rect 12713 20156 13021 20165
rect 12713 20154 12719 20156
rect 12775 20154 12799 20156
rect 12855 20154 12879 20156
rect 12935 20154 12959 20156
rect 13015 20154 13021 20156
rect 12775 20102 12777 20154
rect 12957 20102 12959 20154
rect 12713 20100 12719 20102
rect 12775 20100 12799 20102
rect 12855 20100 12879 20102
rect 12935 20100 12959 20102
rect 13015 20100 13021 20102
rect 12713 20091 13021 20100
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12532 19916 12584 19922
rect 12532 19858 12584 19864
rect 12713 19068 13021 19077
rect 12713 19066 12719 19068
rect 12775 19066 12799 19068
rect 12855 19066 12879 19068
rect 12935 19066 12959 19068
rect 13015 19066 13021 19068
rect 12775 19014 12777 19066
rect 12957 19014 12959 19066
rect 12713 19012 12719 19014
rect 12775 19012 12799 19014
rect 12855 19012 12879 19014
rect 12935 19012 12959 19014
rect 13015 19012 13021 19014
rect 12713 19003 13021 19012
rect 15580 18970 15608 21383
rect 15764 19990 15792 21383
rect 16634 20700 16942 20709
rect 16634 20698 16640 20700
rect 16696 20698 16720 20700
rect 16776 20698 16800 20700
rect 16856 20698 16880 20700
rect 16936 20698 16942 20700
rect 16696 20646 16698 20698
rect 16878 20646 16880 20698
rect 16634 20644 16640 20646
rect 16696 20644 16720 20646
rect 16776 20644 16800 20646
rect 16856 20644 16880 20646
rect 16936 20644 16942 20646
rect 16634 20635 16942 20644
rect 15752 19984 15804 19990
rect 15752 19926 15804 19932
rect 17224 19916 17276 19922
rect 17224 19858 17276 19864
rect 16634 19612 16942 19621
rect 16634 19610 16640 19612
rect 16696 19610 16720 19612
rect 16776 19610 16800 19612
rect 16856 19610 16880 19612
rect 16936 19610 16942 19612
rect 16696 19558 16698 19610
rect 16878 19558 16880 19610
rect 16634 19556 16640 19558
rect 16696 19556 16720 19558
rect 16776 19556 16800 19558
rect 16856 19556 16880 19558
rect 16936 19556 16942 19558
rect 16634 19547 16942 19556
rect 17236 19514 17264 19858
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17512 19242 17540 21383
rect 17866 21312 17922 21321
rect 17922 21270 18000 21298
rect 17866 21247 17922 21256
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 17880 19854 17908 19994
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17500 19236 17552 19242
rect 17500 19178 17552 19184
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 17236 18902 17264 19178
rect 17224 18896 17276 18902
rect 17224 18838 17276 18844
rect 17972 18834 18000 21270
rect 18420 21072 18472 21078
rect 18420 21014 18472 21020
rect 18236 21004 18288 21010
rect 18236 20946 18288 20952
rect 18052 20800 18104 20806
rect 18052 20742 18104 20748
rect 18064 19854 18092 20742
rect 18248 20466 18276 20946
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 18052 19712 18104 19718
rect 18052 19654 18104 19660
rect 18064 19514 18092 19654
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 16634 18524 16942 18533
rect 16634 18522 16640 18524
rect 16696 18522 16720 18524
rect 16776 18522 16800 18524
rect 16856 18522 16880 18524
rect 16936 18522 16942 18524
rect 16696 18470 16698 18522
rect 16878 18470 16880 18522
rect 16634 18468 16640 18470
rect 16696 18468 16720 18470
rect 16776 18468 16800 18470
rect 16856 18468 16880 18470
rect 16936 18468 16942 18470
rect 16634 18459 16942 18468
rect 17052 18358 17080 18702
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 12713 17980 13021 17989
rect 12713 17978 12719 17980
rect 12775 17978 12799 17980
rect 12855 17978 12879 17980
rect 12935 17978 12959 17980
rect 13015 17978 13021 17980
rect 12775 17926 12777 17978
rect 12957 17926 12959 17978
rect 12713 17924 12719 17926
rect 12775 17924 12799 17926
rect 12855 17924 12879 17926
rect 12935 17924 12959 17926
rect 13015 17924 13021 17926
rect 12713 17915 13021 17924
rect 16634 17436 16942 17445
rect 16634 17434 16640 17436
rect 16696 17434 16720 17436
rect 16776 17434 16800 17436
rect 16856 17434 16880 17436
rect 16936 17434 16942 17436
rect 16696 17382 16698 17434
rect 16878 17382 16880 17434
rect 16634 17380 16640 17382
rect 16696 17380 16720 17382
rect 16776 17380 16800 17382
rect 16856 17380 16880 17382
rect 16936 17380 16942 17382
rect 16634 17371 16942 17380
rect 12713 16892 13021 16901
rect 12713 16890 12719 16892
rect 12775 16890 12799 16892
rect 12855 16890 12879 16892
rect 12935 16890 12959 16892
rect 13015 16890 13021 16892
rect 12775 16838 12777 16890
rect 12957 16838 12959 16890
rect 12713 16836 12719 16838
rect 12775 16836 12799 16838
rect 12855 16836 12879 16838
rect 12935 16836 12959 16838
rect 13015 16836 13021 16838
rect 12713 16827 13021 16836
rect 16634 16348 16942 16357
rect 16634 16346 16640 16348
rect 16696 16346 16720 16348
rect 16776 16346 16800 16348
rect 16856 16346 16880 16348
rect 16936 16346 16942 16348
rect 16696 16294 16698 16346
rect 16878 16294 16880 16346
rect 16634 16292 16640 16294
rect 16696 16292 16720 16294
rect 16776 16292 16800 16294
rect 16856 16292 16880 16294
rect 16936 16292 16942 16294
rect 16634 16283 16942 16292
rect 17880 16250 17908 18702
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 18064 15978 18092 19450
rect 18156 16046 18184 20334
rect 18432 20058 18460 21014
rect 19260 20942 19288 21383
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19536 20466 19564 21383
rect 21218 21276 21306 21286
rect 21218 21216 21226 21276
rect 21296 21266 21306 21276
rect 21544 21274 21620 21280
rect 21544 21266 21552 21274
rect 21296 21223 21552 21266
rect 21296 21222 21360 21223
rect 21296 21216 21306 21222
rect 21218 21204 21306 21216
rect 21544 21216 21552 21223
rect 21612 21216 21620 21274
rect 21544 21208 21620 21216
rect 21744 21146 21772 21383
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 19892 21072 19944 21078
rect 19892 21014 19944 21020
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18892 20058 18920 20198
rect 18420 20052 18472 20058
rect 18420 19994 18472 20000
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18432 18766 18460 19994
rect 19248 19848 19300 19854
rect 19300 19796 19564 19802
rect 19248 19790 19564 19796
rect 19260 19786 19564 19790
rect 19812 19786 19840 20810
rect 19904 20330 19932 21014
rect 21088 20936 21140 20942
rect 20902 20904 20958 20913
rect 21088 20878 21140 20884
rect 20902 20839 20958 20848
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20180 20330 20208 20402
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20272 20262 20300 20402
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 20074 20300 20198
rect 19904 20046 20300 20074
rect 19260 19780 19576 19786
rect 19260 19774 19524 19780
rect 19524 19722 19576 19728
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 19536 17202 19564 19722
rect 19904 19514 19932 20046
rect 20364 19854 20392 20402
rect 20555 20156 20863 20165
rect 20555 20154 20561 20156
rect 20617 20154 20641 20156
rect 20697 20154 20721 20156
rect 20777 20154 20801 20156
rect 20857 20154 20863 20156
rect 20617 20102 20619 20154
rect 20799 20102 20801 20154
rect 20555 20100 20561 20102
rect 20617 20100 20641 20102
rect 20697 20100 20721 20102
rect 20777 20100 20801 20102
rect 20857 20100 20863 20102
rect 20555 20091 20863 20100
rect 20812 19984 20864 19990
rect 20810 19952 20812 19961
rect 20864 19952 20866 19961
rect 20810 19887 20866 19896
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19800 19440 19852 19446
rect 19800 19382 19852 19388
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15972 18104 15978
rect 18052 15914 18104 15920
rect 12713 15804 13021 15813
rect 12713 15802 12719 15804
rect 12775 15802 12799 15804
rect 12855 15802 12879 15804
rect 12935 15802 12959 15804
rect 13015 15802 13021 15804
rect 12775 15750 12777 15802
rect 12957 15750 12959 15802
rect 12713 15748 12719 15750
rect 12775 15748 12799 15750
rect 12855 15748 12879 15750
rect 12935 15748 12959 15750
rect 13015 15748 13021 15750
rect 12713 15739 13021 15748
rect 16634 15260 16942 15269
rect 16634 15258 16640 15260
rect 16696 15258 16720 15260
rect 16776 15258 16800 15260
rect 16856 15258 16880 15260
rect 16936 15258 16942 15260
rect 16696 15206 16698 15258
rect 16878 15206 16880 15258
rect 16634 15204 16640 15206
rect 16696 15204 16720 15206
rect 16776 15204 16800 15206
rect 16856 15204 16880 15206
rect 16936 15204 16942 15206
rect 16634 15195 16942 15204
rect 12713 14716 13021 14725
rect 12713 14714 12719 14716
rect 12775 14714 12799 14716
rect 12855 14714 12879 14716
rect 12935 14714 12959 14716
rect 13015 14714 13021 14716
rect 12775 14662 12777 14714
rect 12957 14662 12959 14714
rect 12713 14660 12719 14662
rect 12775 14660 12799 14662
rect 12855 14660 12879 14662
rect 12935 14660 12959 14662
rect 13015 14660 13021 14662
rect 12713 14651 13021 14660
rect 19812 14482 19840 19382
rect 19996 19310 20024 19722
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 20456 14618 20484 19790
rect 20916 19378 20944 20839
rect 20996 20324 21048 20330
rect 20996 20266 21048 20272
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20628 19304 20680 19310
rect 20626 19272 20628 19281
rect 20680 19272 20682 19281
rect 20626 19207 20682 19216
rect 20555 19068 20863 19077
rect 20555 19066 20561 19068
rect 20617 19066 20641 19068
rect 20697 19066 20721 19068
rect 20777 19066 20801 19068
rect 20857 19066 20863 19068
rect 20617 19014 20619 19066
rect 20799 19014 20801 19066
rect 20555 19012 20561 19014
rect 20617 19012 20641 19014
rect 20697 19012 20721 19014
rect 20777 19012 20801 19014
rect 20857 19012 20863 19014
rect 20555 19003 20863 19012
rect 20555 17980 20863 17989
rect 20555 17978 20561 17980
rect 20617 17978 20641 17980
rect 20697 17978 20721 17980
rect 20777 17978 20801 17980
rect 20857 17978 20863 17980
rect 20617 17926 20619 17978
rect 20799 17926 20801 17978
rect 20555 17924 20561 17926
rect 20617 17924 20641 17926
rect 20697 17924 20721 17926
rect 20777 17924 20801 17926
rect 20857 17924 20863 17926
rect 20555 17915 20863 17924
rect 20555 16892 20863 16901
rect 20555 16890 20561 16892
rect 20617 16890 20641 16892
rect 20697 16890 20721 16892
rect 20777 16890 20801 16892
rect 20857 16890 20863 16892
rect 20617 16838 20619 16890
rect 20799 16838 20801 16890
rect 20555 16836 20561 16838
rect 20617 16836 20641 16838
rect 20697 16836 20721 16838
rect 20777 16836 20801 16838
rect 20857 16836 20863 16838
rect 20555 16827 20863 16836
rect 21008 16114 21036 20266
rect 21100 19990 21128 20878
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21088 19984 21140 19990
rect 21192 19961 21220 20334
rect 21088 19926 21140 19932
rect 21178 19952 21234 19961
rect 21178 19887 21234 19896
rect 21548 19848 21600 19854
rect 21548 19790 21600 19796
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21468 19174 21496 19246
rect 21456 19168 21508 19174
rect 21456 19110 21508 19116
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20555 15804 20863 15813
rect 20555 15802 20561 15804
rect 20617 15802 20641 15804
rect 20697 15802 20721 15804
rect 20777 15802 20801 15804
rect 20857 15802 20863 15804
rect 20617 15750 20619 15802
rect 20799 15750 20801 15802
rect 20555 15748 20561 15750
rect 20617 15748 20641 15750
rect 20697 15748 20721 15750
rect 20777 15748 20801 15750
rect 20857 15748 20863 15750
rect 20555 15739 20863 15748
rect 20555 14716 20863 14725
rect 20555 14714 20561 14716
rect 20617 14714 20641 14716
rect 20697 14714 20721 14716
rect 20777 14714 20801 14716
rect 20857 14714 20863 14716
rect 20617 14662 20619 14714
rect 20799 14662 20801 14714
rect 20555 14660 20561 14662
rect 20617 14660 20641 14662
rect 20697 14660 20721 14662
rect 20777 14660 20801 14662
rect 20857 14660 20863 14662
rect 20555 14651 20863 14660
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 19800 14476 19852 14482
rect 19800 14418 19852 14424
rect 20168 14476 20220 14482
rect 20168 14418 20220 14424
rect 16634 14172 16942 14181
rect 16634 14170 16640 14172
rect 16696 14170 16720 14172
rect 16776 14170 16800 14172
rect 16856 14170 16880 14172
rect 16936 14170 16942 14172
rect 16696 14118 16698 14170
rect 16878 14118 16880 14170
rect 16634 14116 16640 14118
rect 16696 14116 16720 14118
rect 16776 14116 16800 14118
rect 16856 14116 16880 14118
rect 16936 14116 16942 14118
rect 16634 14107 16942 14116
rect 20180 14006 20208 14418
rect 20168 14000 20220 14006
rect 20168 13942 20220 13948
rect 12713 13628 13021 13637
rect 12713 13626 12719 13628
rect 12775 13626 12799 13628
rect 12855 13626 12879 13628
rect 12935 13626 12959 13628
rect 13015 13626 13021 13628
rect 12775 13574 12777 13626
rect 12957 13574 12959 13626
rect 12713 13572 12719 13574
rect 12775 13572 12799 13574
rect 12855 13572 12879 13574
rect 12935 13572 12959 13574
rect 13015 13572 13021 13574
rect 12713 13563 13021 13572
rect 16634 13084 16942 13093
rect 16634 13082 16640 13084
rect 16696 13082 16720 13084
rect 16776 13082 16800 13084
rect 16856 13082 16880 13084
rect 16936 13082 16942 13084
rect 16696 13030 16698 13082
rect 16878 13030 16880 13082
rect 16634 13028 16640 13030
rect 16696 13028 16720 13030
rect 16776 13028 16800 13030
rect 16856 13028 16880 13030
rect 16936 13028 16942 13030
rect 16634 13019 16942 13028
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 4871 12540 5179 12549
rect 4871 12538 4877 12540
rect 4933 12538 4957 12540
rect 5013 12538 5037 12540
rect 5093 12538 5117 12540
rect 5173 12538 5179 12540
rect 4933 12486 4935 12538
rect 5115 12486 5117 12538
rect 4871 12484 4877 12486
rect 4933 12484 4957 12486
rect 5013 12484 5037 12486
rect 5093 12484 5117 12486
rect 5173 12484 5179 12486
rect 4871 12475 5179 12484
rect 12713 12540 13021 12549
rect 12713 12538 12719 12540
rect 12775 12538 12799 12540
rect 12855 12538 12879 12540
rect 12935 12538 12959 12540
rect 13015 12538 13021 12540
rect 12775 12486 12777 12538
rect 12957 12486 12959 12538
rect 12713 12484 12719 12486
rect 12775 12484 12799 12486
rect 12855 12484 12879 12486
rect 12935 12484 12959 12486
rect 13015 12484 13021 12486
rect 12713 12475 13021 12484
rect 20180 12170 20208 13942
rect 20555 13628 20863 13637
rect 20555 13626 20561 13628
rect 20617 13626 20641 13628
rect 20697 13626 20721 13628
rect 20777 13626 20801 13628
rect 20857 13626 20863 13628
rect 20617 13574 20619 13626
rect 20799 13574 20801 13626
rect 20555 13572 20561 13574
rect 20617 13572 20641 13574
rect 20697 13572 20721 13574
rect 20777 13572 20801 13574
rect 20857 13572 20863 13574
rect 20555 13563 20863 13572
rect 20555 12540 20863 12549
rect 20555 12538 20561 12540
rect 20617 12538 20641 12540
rect 20697 12538 20721 12540
rect 20777 12538 20801 12540
rect 20857 12538 20863 12540
rect 20617 12486 20619 12538
rect 20799 12486 20801 12538
rect 20555 12484 20561 12486
rect 20617 12484 20641 12486
rect 20697 12484 20721 12486
rect 20777 12484 20801 12486
rect 20857 12484 20863 12486
rect 20555 12475 20863 12484
rect 21008 12442 21036 16050
rect 21560 15162 21588 19790
rect 21640 19712 21692 19718
rect 21640 19654 21692 19660
rect 21652 19310 21680 19654
rect 21836 19553 21864 19790
rect 21822 19544 21878 19553
rect 21822 19479 21878 19488
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21928 18698 21956 20334
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22020 19281 22048 19450
rect 22006 19272 22062 19281
rect 22006 19207 22062 19216
rect 22112 18766 22140 19450
rect 22204 19242 22232 20742
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 22296 19922 22324 20538
rect 22376 20460 22428 20466
rect 22376 20402 22428 20408
rect 22284 19916 22336 19922
rect 22284 19858 22336 19864
rect 22192 19236 22244 19242
rect 22192 19178 22244 19184
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 18766 22324 19110
rect 22100 18760 22152 18766
rect 22100 18702 22152 18708
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 22388 17202 22416 20402
rect 22480 19378 22508 20810
rect 22652 20528 22704 20534
rect 22652 20470 22704 20476
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22664 17882 22692 20470
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22756 19514 22784 20334
rect 22836 19984 22888 19990
rect 22836 19926 22888 19932
rect 22848 19854 22876 19926
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22756 18970 22784 19246
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22940 18766 22968 21383
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23020 19508 23072 19514
rect 23020 19450 23072 19456
rect 23032 19174 23060 19450
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 23124 18834 23152 20946
rect 23676 20534 23704 21383
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23756 20596 23808 20602
rect 23756 20538 23808 20544
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23400 20058 23428 20334
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23308 19446 23336 19654
rect 23296 19440 23348 19446
rect 23296 19382 23348 19388
rect 23400 19378 23428 19994
rect 23492 19990 23520 20266
rect 23480 19984 23532 19990
rect 23480 19926 23532 19932
rect 23584 19786 23612 20402
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23570 19544 23626 19553
rect 23570 19479 23626 19488
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 19304 23348 19310
rect 23348 19252 23520 19258
rect 23296 19246 23520 19252
rect 23308 19230 23520 19246
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 22928 18760 22980 18766
rect 22928 18702 22980 18708
rect 22652 17876 22704 17882
rect 22652 17818 22704 17824
rect 22664 17202 22692 17818
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 22388 16794 22416 17138
rect 23124 17134 23152 18770
rect 23492 18766 23520 19230
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23480 18624 23532 18630
rect 23480 18566 23532 18572
rect 23492 17882 23520 18566
rect 23584 18426 23612 19479
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23572 17740 23624 17746
rect 23572 17682 23624 17688
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 23584 16522 23612 17682
rect 23676 17338 23704 19382
rect 23768 19310 23796 20538
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23756 18760 23808 18766
rect 23756 18702 23808 18708
rect 23664 17332 23716 17338
rect 23664 17274 23716 17280
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 20996 12436 21048 12442
rect 21560 12434 21588 15098
rect 23676 14958 23704 17274
rect 23664 14952 23716 14958
rect 23664 14894 23716 14900
rect 23768 12850 23796 18702
rect 23860 17678 23888 20538
rect 24044 20466 24072 21082
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 23952 17746 23980 19926
rect 24136 19258 24164 21014
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24228 19378 24256 20402
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24136 19242 24256 19258
rect 24136 19236 24268 19242
rect 24136 19230 24216 19236
rect 24032 18284 24084 18290
rect 24032 18226 24084 18232
rect 23940 17740 23992 17746
rect 23940 17682 23992 17688
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 23860 16590 23888 17614
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23952 15094 23980 17138
rect 24044 16454 24072 18226
rect 24136 17202 24164 19230
rect 24216 19178 24268 19184
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 24124 17196 24176 17202
rect 24124 17138 24176 17144
rect 24124 16516 24176 16522
rect 24124 16458 24176 16464
rect 24032 16448 24084 16454
rect 24032 16390 24084 16396
rect 23940 15088 23992 15094
rect 23940 15030 23992 15036
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 21640 12436 21692 12442
rect 21560 12406 21640 12434
rect 20996 12378 21048 12384
rect 21640 12378 21692 12384
rect 24044 12306 24072 16390
rect 24136 15026 24164 16458
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24228 12646 24256 18634
rect 24320 16658 24348 20538
rect 24412 19922 24440 21383
rect 24476 20700 24784 20709
rect 24476 20698 24482 20700
rect 24538 20698 24562 20700
rect 24618 20698 24642 20700
rect 24698 20698 24722 20700
rect 24778 20698 24784 20700
rect 24538 20646 24540 20698
rect 24720 20646 24722 20698
rect 24476 20644 24482 20646
rect 24538 20644 24562 20646
rect 24618 20644 24642 20646
rect 24698 20644 24722 20646
rect 24778 20644 24784 20646
rect 24476 20635 24784 20644
rect 24766 20496 24822 20505
rect 25884 20466 25912 21383
rect 27342 21040 27398 21049
rect 27342 20975 27398 20984
rect 27356 20466 27384 20975
rect 27448 20466 27476 21383
rect 28630 21040 28686 21049
rect 28630 20975 28686 20984
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28460 20602 28488 20810
rect 28448 20596 28500 20602
rect 28448 20538 28500 20544
rect 28644 20466 28672 20975
rect 24766 20431 24822 20440
rect 25872 20460 25924 20466
rect 24492 20392 24544 20398
rect 24492 20334 24544 20340
rect 24400 19916 24452 19922
rect 24400 19858 24452 19864
rect 24504 19700 24532 20334
rect 24780 19854 24808 20431
rect 25872 20402 25924 20408
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27436 20460 27488 20466
rect 27436 20402 27488 20408
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 25136 20256 25188 20262
rect 25136 20198 25188 20204
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24412 19672 24532 19700
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 24320 15042 24348 16594
rect 24412 16522 24440 19672
rect 24476 19612 24784 19621
rect 24476 19610 24482 19612
rect 24538 19610 24562 19612
rect 24618 19610 24642 19612
rect 24698 19610 24722 19612
rect 24778 19610 24784 19612
rect 24538 19558 24540 19610
rect 24720 19558 24722 19610
rect 24476 19556 24482 19558
rect 24538 19556 24562 19558
rect 24618 19556 24642 19558
rect 24698 19556 24722 19558
rect 24778 19556 24784 19558
rect 24476 19547 24784 19556
rect 24872 19378 24900 20198
rect 24860 19372 24912 19378
rect 24860 19314 24912 19320
rect 24476 18524 24784 18533
rect 24476 18522 24482 18524
rect 24538 18522 24562 18524
rect 24618 18522 24642 18524
rect 24698 18522 24722 18524
rect 24778 18522 24784 18524
rect 24538 18470 24540 18522
rect 24720 18470 24722 18522
rect 24476 18468 24482 18470
rect 24538 18468 24562 18470
rect 24618 18468 24642 18470
rect 24698 18468 24722 18470
rect 24778 18468 24784 18470
rect 24476 18459 24784 18468
rect 24476 17436 24784 17445
rect 24476 17434 24482 17436
rect 24538 17434 24562 17436
rect 24618 17434 24642 17436
rect 24698 17434 24722 17436
rect 24778 17434 24784 17436
rect 24538 17382 24540 17434
rect 24720 17382 24722 17434
rect 24476 17380 24482 17382
rect 24538 17380 24562 17382
rect 24618 17380 24642 17382
rect 24698 17380 24722 17382
rect 24778 17380 24784 17382
rect 24476 17371 24784 17380
rect 25148 17270 25176 20198
rect 25412 19712 25464 19718
rect 25412 19654 25464 19660
rect 25320 18352 25372 18358
rect 25320 18294 25372 18300
rect 25136 17264 25188 17270
rect 25136 17206 25188 17212
rect 24400 16516 24452 16522
rect 24400 16458 24452 16464
rect 24476 16348 24784 16357
rect 24476 16346 24482 16348
rect 24538 16346 24562 16348
rect 24618 16346 24642 16348
rect 24698 16346 24722 16348
rect 24778 16346 24784 16348
rect 24538 16294 24540 16346
rect 24720 16294 24722 16346
rect 24476 16292 24482 16294
rect 24538 16292 24562 16294
rect 24618 16292 24642 16294
rect 24698 16292 24722 16294
rect 24778 16292 24784 16294
rect 24476 16283 24784 16292
rect 24476 15260 24784 15269
rect 24476 15258 24482 15260
rect 24538 15258 24562 15260
rect 24618 15258 24642 15260
rect 24698 15258 24722 15260
rect 24778 15258 24784 15260
rect 24538 15206 24540 15258
rect 24720 15206 24722 15258
rect 24476 15204 24482 15206
rect 24538 15204 24562 15206
rect 24618 15204 24642 15206
rect 24698 15204 24722 15206
rect 24778 15204 24784 15206
rect 24476 15195 24784 15204
rect 24320 15026 24440 15042
rect 25148 15026 25176 17206
rect 25332 15162 25360 18294
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 24320 15020 24452 15026
rect 24320 15014 24400 15020
rect 24400 14962 24452 14968
rect 25136 15020 25188 15026
rect 25136 14962 25188 14968
rect 24476 14172 24784 14181
rect 24476 14170 24482 14172
rect 24538 14170 24562 14172
rect 24618 14170 24642 14172
rect 24698 14170 24722 14172
rect 24778 14170 24784 14172
rect 24538 14118 24540 14170
rect 24720 14118 24722 14170
rect 24476 14116 24482 14118
rect 24538 14116 24562 14118
rect 24618 14116 24642 14118
rect 24698 14116 24722 14118
rect 24778 14116 24784 14118
rect 24476 14107 24784 14116
rect 25424 14006 25452 19654
rect 27172 19514 27200 20198
rect 27816 19990 27844 20198
rect 28397 20156 28705 20165
rect 28397 20154 28403 20156
rect 28459 20154 28483 20156
rect 28539 20154 28563 20156
rect 28619 20154 28643 20156
rect 28699 20154 28705 20156
rect 28459 20102 28461 20154
rect 28641 20102 28643 20154
rect 28397 20100 28403 20102
rect 28459 20100 28483 20102
rect 28539 20100 28563 20102
rect 28619 20100 28643 20102
rect 28699 20100 28705 20102
rect 28397 20091 28705 20100
rect 27804 19984 27856 19990
rect 27804 19926 27856 19932
rect 28828 19854 28856 21383
rect 29918 21040 29974 21049
rect 29918 20975 29974 20984
rect 29932 20466 29960 20975
rect 30300 20466 30328 21383
rect 33598 21280 33714 21294
rect 33598 21208 33614 21280
rect 33696 21208 33714 21280
rect 33598 21192 33714 21208
rect 32318 20700 32626 20709
rect 32318 20698 32324 20700
rect 32380 20698 32404 20700
rect 32460 20698 32484 20700
rect 32540 20698 32564 20700
rect 32620 20698 32626 20700
rect 32380 20646 32382 20698
rect 32562 20646 32564 20698
rect 32318 20644 32324 20646
rect 32380 20644 32404 20646
rect 32460 20644 32484 20646
rect 32540 20644 32564 20646
rect 32620 20644 32626 20646
rect 32318 20635 32626 20644
rect 29920 20460 29972 20466
rect 29920 20402 29972 20408
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 27160 19508 27212 19514
rect 27160 19450 27212 19456
rect 28397 19068 28705 19077
rect 28397 19066 28403 19068
rect 28459 19066 28483 19068
rect 28539 19066 28563 19068
rect 28619 19066 28643 19068
rect 28699 19066 28705 19068
rect 28459 19014 28461 19066
rect 28641 19014 28643 19066
rect 28397 19012 28403 19014
rect 28459 19012 28483 19014
rect 28539 19012 28563 19014
rect 28619 19012 28643 19014
rect 28699 19012 28705 19014
rect 28397 19003 28705 19012
rect 28397 17980 28705 17989
rect 28397 17978 28403 17980
rect 28459 17978 28483 17980
rect 28539 17978 28563 17980
rect 28619 17978 28643 17980
rect 28699 17978 28705 17980
rect 28459 17926 28461 17978
rect 28641 17926 28643 17978
rect 28397 17924 28403 17926
rect 28459 17924 28483 17926
rect 28539 17924 28563 17926
rect 28619 17924 28643 17926
rect 28699 17924 28705 17926
rect 28397 17915 28705 17924
rect 28397 16892 28705 16901
rect 28397 16890 28403 16892
rect 28459 16890 28483 16892
rect 28539 16890 28563 16892
rect 28619 16890 28643 16892
rect 28699 16890 28705 16892
rect 28459 16838 28461 16890
rect 28641 16838 28643 16890
rect 28397 16836 28403 16838
rect 28459 16836 28483 16838
rect 28539 16836 28563 16838
rect 28619 16836 28643 16838
rect 28699 16836 28705 16838
rect 28397 16827 28705 16836
rect 28397 15804 28705 15813
rect 28397 15802 28403 15804
rect 28459 15802 28483 15804
rect 28539 15802 28563 15804
rect 28619 15802 28643 15804
rect 28699 15802 28705 15804
rect 28459 15750 28461 15802
rect 28641 15750 28643 15802
rect 28397 15748 28403 15750
rect 28459 15748 28483 15750
rect 28539 15748 28563 15750
rect 28619 15748 28643 15750
rect 28699 15748 28705 15750
rect 28397 15739 28705 15748
rect 28397 14716 28705 14725
rect 28397 14714 28403 14716
rect 28459 14714 28483 14716
rect 28539 14714 28563 14716
rect 28619 14714 28643 14716
rect 28699 14714 28705 14716
rect 28459 14662 28461 14714
rect 28641 14662 28643 14714
rect 28397 14660 28403 14662
rect 28459 14660 28483 14662
rect 28539 14660 28563 14662
rect 28619 14660 28643 14662
rect 28699 14660 28705 14662
rect 28397 14651 28705 14660
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25516 14074 25544 14350
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 30392 14006 30420 20198
rect 32318 19612 32626 19621
rect 32318 19610 32324 19612
rect 32380 19610 32404 19612
rect 32460 19610 32484 19612
rect 32540 19610 32564 19612
rect 32620 19610 32626 19612
rect 32380 19558 32382 19610
rect 32562 19558 32564 19610
rect 32318 19556 32324 19558
rect 32380 19556 32404 19558
rect 32460 19556 32484 19558
rect 32540 19556 32564 19558
rect 32620 19556 32626 19558
rect 32318 19547 32626 19556
rect 32318 18524 32626 18533
rect 32318 18522 32324 18524
rect 32380 18522 32404 18524
rect 32460 18522 32484 18524
rect 32540 18522 32564 18524
rect 32620 18522 32626 18524
rect 32380 18470 32382 18522
rect 32562 18470 32564 18522
rect 32318 18468 32324 18470
rect 32380 18468 32404 18470
rect 32460 18468 32484 18470
rect 32540 18468 32564 18470
rect 32620 18468 32626 18470
rect 32318 18459 32626 18468
rect 32318 17436 32626 17445
rect 32318 17434 32324 17436
rect 32380 17434 32404 17436
rect 32460 17434 32484 17436
rect 32540 17434 32564 17436
rect 32620 17434 32626 17436
rect 32380 17382 32382 17434
rect 32562 17382 32564 17434
rect 32318 17380 32324 17382
rect 32380 17380 32404 17382
rect 32460 17380 32484 17382
rect 32540 17380 32564 17382
rect 32620 17380 32626 17382
rect 32318 17371 32626 17380
rect 32318 16348 32626 16357
rect 32318 16346 32324 16348
rect 32380 16346 32404 16348
rect 32460 16346 32484 16348
rect 32540 16346 32564 16348
rect 32620 16346 32626 16348
rect 32380 16294 32382 16346
rect 32562 16294 32564 16346
rect 32318 16292 32324 16294
rect 32380 16292 32404 16294
rect 32460 16292 32484 16294
rect 32540 16292 32564 16294
rect 32620 16292 32626 16294
rect 32318 16283 32626 16292
rect 32318 15260 32626 15269
rect 32318 15258 32324 15260
rect 32380 15258 32404 15260
rect 32460 15258 32484 15260
rect 32540 15258 32564 15260
rect 32620 15258 32626 15260
rect 32380 15206 32382 15258
rect 32562 15206 32564 15258
rect 32318 15204 32324 15206
rect 32380 15204 32404 15206
rect 32460 15204 32484 15206
rect 32540 15204 32564 15206
rect 32620 15204 32626 15206
rect 32318 15195 32626 15204
rect 32318 14172 32626 14181
rect 32318 14170 32324 14172
rect 32380 14170 32404 14172
rect 32460 14170 32484 14172
rect 32540 14170 32564 14172
rect 32620 14170 32626 14172
rect 32380 14118 32382 14170
rect 32562 14118 32564 14170
rect 32318 14116 32324 14118
rect 32380 14116 32404 14118
rect 32460 14116 32484 14118
rect 32540 14116 32564 14118
rect 32620 14116 32626 14118
rect 32318 14107 32626 14116
rect 25412 14000 25464 14006
rect 25412 13942 25464 13948
rect 30380 14000 30432 14006
rect 30380 13942 30432 13948
rect 28397 13628 28705 13637
rect 28397 13626 28403 13628
rect 28459 13626 28483 13628
rect 28539 13626 28563 13628
rect 28619 13626 28643 13628
rect 28699 13626 28705 13628
rect 28459 13574 28461 13626
rect 28641 13574 28643 13626
rect 28397 13572 28403 13574
rect 28459 13572 28483 13574
rect 28539 13572 28563 13574
rect 28619 13572 28643 13574
rect 28699 13572 28705 13574
rect 28397 13563 28705 13572
rect 24476 13084 24784 13093
rect 24476 13082 24482 13084
rect 24538 13082 24562 13084
rect 24618 13082 24642 13084
rect 24698 13082 24722 13084
rect 24778 13082 24784 13084
rect 24538 13030 24540 13082
rect 24720 13030 24722 13082
rect 24476 13028 24482 13030
rect 24538 13028 24562 13030
rect 24618 13028 24642 13030
rect 24698 13028 24722 13030
rect 24778 13028 24784 13030
rect 24476 13019 24784 13028
rect 32318 13084 32626 13093
rect 32318 13082 32324 13084
rect 32380 13082 32404 13084
rect 32460 13082 32484 13084
rect 32540 13082 32564 13084
rect 32620 13082 32626 13084
rect 32380 13030 32382 13082
rect 32562 13030 32564 13082
rect 32318 13028 32324 13030
rect 32380 13028 32404 13030
rect 32460 13028 32484 13030
rect 32540 13028 32564 13030
rect 32620 13028 32626 13030
rect 32318 13019 32626 13028
rect 24216 12640 24268 12646
rect 24216 12582 24268 12588
rect 28397 12540 28705 12549
rect 28397 12538 28403 12540
rect 28459 12538 28483 12540
rect 28539 12538 28563 12540
rect 28619 12538 28643 12540
rect 28699 12538 28705 12540
rect 28459 12486 28461 12538
rect 28641 12486 28643 12538
rect 28397 12484 28403 12486
rect 28459 12484 28483 12486
rect 28539 12484 28563 12486
rect 28619 12484 28643 12486
rect 28699 12484 28705 12486
rect 28397 12475 28705 12484
rect 24032 12300 24084 12306
rect 24032 12242 24084 12248
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 8792 11996 9100 12005
rect 8792 11994 8798 11996
rect 8854 11994 8878 11996
rect 8934 11994 8958 11996
rect 9014 11994 9038 11996
rect 9094 11994 9100 11996
rect 8854 11942 8856 11994
rect 9036 11942 9038 11994
rect 8792 11940 8798 11942
rect 8854 11940 8878 11942
rect 8934 11940 8958 11942
rect 9014 11940 9038 11942
rect 9094 11940 9100 11942
rect 8792 11931 9100 11940
rect 16634 11996 16942 12005
rect 16634 11994 16640 11996
rect 16696 11994 16720 11996
rect 16776 11994 16800 11996
rect 16856 11994 16880 11996
rect 16936 11994 16942 11996
rect 16696 11942 16698 11994
rect 16878 11942 16880 11994
rect 16634 11940 16640 11942
rect 16696 11940 16720 11942
rect 16776 11940 16800 11942
rect 16856 11940 16880 11942
rect 16936 11940 16942 11942
rect 16634 11931 16942 11940
rect 24476 11996 24784 12005
rect 24476 11994 24482 11996
rect 24538 11994 24562 11996
rect 24618 11994 24642 11996
rect 24698 11994 24722 11996
rect 24778 11994 24784 11996
rect 24538 11942 24540 11994
rect 24720 11942 24722 11994
rect 24476 11940 24482 11942
rect 24538 11940 24562 11942
rect 24618 11940 24642 11942
rect 24698 11940 24722 11942
rect 24778 11940 24784 11942
rect 24476 11931 24784 11940
rect 32318 11996 32626 12005
rect 32318 11994 32324 11996
rect 32380 11994 32404 11996
rect 32460 11994 32484 11996
rect 32540 11994 32564 11996
rect 32620 11994 32626 11996
rect 32380 11942 32382 11994
rect 32562 11942 32564 11994
rect 32318 11940 32324 11942
rect 32380 11940 32404 11942
rect 32460 11940 32484 11942
rect 32540 11940 32564 11942
rect 32620 11940 32626 11942
rect 32318 11931 32626 11940
rect 4871 11452 5179 11461
rect 4871 11450 4877 11452
rect 4933 11450 4957 11452
rect 5013 11450 5037 11452
rect 5093 11450 5117 11452
rect 5173 11450 5179 11452
rect 4933 11398 4935 11450
rect 5115 11398 5117 11450
rect 4871 11396 4877 11398
rect 4933 11396 4957 11398
rect 5013 11396 5037 11398
rect 5093 11396 5117 11398
rect 5173 11396 5179 11398
rect 4871 11387 5179 11396
rect 12713 11452 13021 11461
rect 12713 11450 12719 11452
rect 12775 11450 12799 11452
rect 12855 11450 12879 11452
rect 12935 11450 12959 11452
rect 13015 11450 13021 11452
rect 12775 11398 12777 11450
rect 12957 11398 12959 11450
rect 12713 11396 12719 11398
rect 12775 11396 12799 11398
rect 12855 11396 12879 11398
rect 12935 11396 12959 11398
rect 13015 11396 13021 11398
rect 12713 11387 13021 11396
rect 20555 11452 20863 11461
rect 20555 11450 20561 11452
rect 20617 11450 20641 11452
rect 20697 11450 20721 11452
rect 20777 11450 20801 11452
rect 20857 11450 20863 11452
rect 20617 11398 20619 11450
rect 20799 11398 20801 11450
rect 20555 11396 20561 11398
rect 20617 11396 20641 11398
rect 20697 11396 20721 11398
rect 20777 11396 20801 11398
rect 20857 11396 20863 11398
rect 20555 11387 20863 11396
rect 28397 11452 28705 11461
rect 28397 11450 28403 11452
rect 28459 11450 28483 11452
rect 28539 11450 28563 11452
rect 28619 11450 28643 11452
rect 28699 11450 28705 11452
rect 28459 11398 28461 11450
rect 28641 11398 28643 11450
rect 28397 11396 28403 11398
rect 28459 11396 28483 11398
rect 28539 11396 28563 11398
rect 28619 11396 28643 11398
rect 28699 11396 28705 11398
rect 28397 11387 28705 11396
rect 8792 10908 9100 10917
rect 8792 10906 8798 10908
rect 8854 10906 8878 10908
rect 8934 10906 8958 10908
rect 9014 10906 9038 10908
rect 9094 10906 9100 10908
rect 8854 10854 8856 10906
rect 9036 10854 9038 10906
rect 8792 10852 8798 10854
rect 8854 10852 8878 10854
rect 8934 10852 8958 10854
rect 9014 10852 9038 10854
rect 9094 10852 9100 10854
rect 8792 10843 9100 10852
rect 16634 10908 16942 10917
rect 16634 10906 16640 10908
rect 16696 10906 16720 10908
rect 16776 10906 16800 10908
rect 16856 10906 16880 10908
rect 16936 10906 16942 10908
rect 16696 10854 16698 10906
rect 16878 10854 16880 10906
rect 16634 10852 16640 10854
rect 16696 10852 16720 10854
rect 16776 10852 16800 10854
rect 16856 10852 16880 10854
rect 16936 10852 16942 10854
rect 16634 10843 16942 10852
rect 24476 10908 24784 10917
rect 24476 10906 24482 10908
rect 24538 10906 24562 10908
rect 24618 10906 24642 10908
rect 24698 10906 24722 10908
rect 24778 10906 24784 10908
rect 24538 10854 24540 10906
rect 24720 10854 24722 10906
rect 24476 10852 24482 10854
rect 24538 10852 24562 10854
rect 24618 10852 24642 10854
rect 24698 10852 24722 10854
rect 24778 10852 24784 10854
rect 24476 10843 24784 10852
rect 32318 10908 32626 10917
rect 32318 10906 32324 10908
rect 32380 10906 32404 10908
rect 32460 10906 32484 10908
rect 32540 10906 32564 10908
rect 32620 10906 32626 10908
rect 32380 10854 32382 10906
rect 32562 10854 32564 10906
rect 32318 10852 32324 10854
rect 32380 10852 32404 10854
rect 32460 10852 32484 10854
rect 32540 10852 32564 10854
rect 32620 10852 32626 10854
rect 32318 10843 32626 10852
rect 4871 10364 5179 10373
rect 4871 10362 4877 10364
rect 4933 10362 4957 10364
rect 5013 10362 5037 10364
rect 5093 10362 5117 10364
rect 5173 10362 5179 10364
rect 4933 10310 4935 10362
rect 5115 10310 5117 10362
rect 4871 10308 4877 10310
rect 4933 10308 4957 10310
rect 5013 10308 5037 10310
rect 5093 10308 5117 10310
rect 5173 10308 5179 10310
rect 4871 10299 5179 10308
rect 12713 10364 13021 10373
rect 12713 10362 12719 10364
rect 12775 10362 12799 10364
rect 12855 10362 12879 10364
rect 12935 10362 12959 10364
rect 13015 10362 13021 10364
rect 12775 10310 12777 10362
rect 12957 10310 12959 10362
rect 12713 10308 12719 10310
rect 12775 10308 12799 10310
rect 12855 10308 12879 10310
rect 12935 10308 12959 10310
rect 13015 10308 13021 10310
rect 12713 10299 13021 10308
rect 20555 10364 20863 10373
rect 20555 10362 20561 10364
rect 20617 10362 20641 10364
rect 20697 10362 20721 10364
rect 20777 10362 20801 10364
rect 20857 10362 20863 10364
rect 20617 10310 20619 10362
rect 20799 10310 20801 10362
rect 20555 10308 20561 10310
rect 20617 10308 20641 10310
rect 20697 10308 20721 10310
rect 20777 10308 20801 10310
rect 20857 10308 20863 10310
rect 20555 10299 20863 10308
rect 28397 10364 28705 10373
rect 28397 10362 28403 10364
rect 28459 10362 28483 10364
rect 28539 10362 28563 10364
rect 28619 10362 28643 10364
rect 28699 10362 28705 10364
rect 28459 10310 28461 10362
rect 28641 10310 28643 10362
rect 28397 10308 28403 10310
rect 28459 10308 28483 10310
rect 28539 10308 28563 10310
rect 28619 10308 28643 10310
rect 28699 10308 28705 10310
rect 28397 10299 28705 10308
rect 8792 9820 9100 9829
rect 8792 9818 8798 9820
rect 8854 9818 8878 9820
rect 8934 9818 8958 9820
rect 9014 9818 9038 9820
rect 9094 9818 9100 9820
rect 8854 9766 8856 9818
rect 9036 9766 9038 9818
rect 8792 9764 8798 9766
rect 8854 9764 8878 9766
rect 8934 9764 8958 9766
rect 9014 9764 9038 9766
rect 9094 9764 9100 9766
rect 8792 9755 9100 9764
rect 16634 9820 16942 9829
rect 16634 9818 16640 9820
rect 16696 9818 16720 9820
rect 16776 9818 16800 9820
rect 16856 9818 16880 9820
rect 16936 9818 16942 9820
rect 16696 9766 16698 9818
rect 16878 9766 16880 9818
rect 16634 9764 16640 9766
rect 16696 9764 16720 9766
rect 16776 9764 16800 9766
rect 16856 9764 16880 9766
rect 16936 9764 16942 9766
rect 16634 9755 16942 9764
rect 24476 9820 24784 9829
rect 24476 9818 24482 9820
rect 24538 9818 24562 9820
rect 24618 9818 24642 9820
rect 24698 9818 24722 9820
rect 24778 9818 24784 9820
rect 24538 9766 24540 9818
rect 24720 9766 24722 9818
rect 24476 9764 24482 9766
rect 24538 9764 24562 9766
rect 24618 9764 24642 9766
rect 24698 9764 24722 9766
rect 24778 9764 24784 9766
rect 24476 9755 24784 9764
rect 32318 9820 32626 9829
rect 32318 9818 32324 9820
rect 32380 9818 32404 9820
rect 32460 9818 32484 9820
rect 32540 9818 32564 9820
rect 32620 9818 32626 9820
rect 32380 9766 32382 9818
rect 32562 9766 32564 9818
rect 32318 9764 32324 9766
rect 32380 9764 32404 9766
rect 32460 9764 32484 9766
rect 32540 9764 32564 9766
rect 32620 9764 32626 9766
rect 32318 9755 32626 9764
rect 4871 9276 5179 9285
rect 4871 9274 4877 9276
rect 4933 9274 4957 9276
rect 5013 9274 5037 9276
rect 5093 9274 5117 9276
rect 5173 9274 5179 9276
rect 4933 9222 4935 9274
rect 5115 9222 5117 9274
rect 4871 9220 4877 9222
rect 4933 9220 4957 9222
rect 5013 9220 5037 9222
rect 5093 9220 5117 9222
rect 5173 9220 5179 9222
rect 4871 9211 5179 9220
rect 12713 9276 13021 9285
rect 12713 9274 12719 9276
rect 12775 9274 12799 9276
rect 12855 9274 12879 9276
rect 12935 9274 12959 9276
rect 13015 9274 13021 9276
rect 12775 9222 12777 9274
rect 12957 9222 12959 9274
rect 12713 9220 12719 9222
rect 12775 9220 12799 9222
rect 12855 9220 12879 9222
rect 12935 9220 12959 9222
rect 13015 9220 13021 9222
rect 12713 9211 13021 9220
rect 20555 9276 20863 9285
rect 20555 9274 20561 9276
rect 20617 9274 20641 9276
rect 20697 9274 20721 9276
rect 20777 9274 20801 9276
rect 20857 9274 20863 9276
rect 20617 9222 20619 9274
rect 20799 9222 20801 9274
rect 20555 9220 20561 9222
rect 20617 9220 20641 9222
rect 20697 9220 20721 9222
rect 20777 9220 20801 9222
rect 20857 9220 20863 9222
rect 20555 9211 20863 9220
rect 28397 9276 28705 9285
rect 28397 9274 28403 9276
rect 28459 9274 28483 9276
rect 28539 9274 28563 9276
rect 28619 9274 28643 9276
rect 28699 9274 28705 9276
rect 28459 9222 28461 9274
rect 28641 9222 28643 9274
rect 28397 9220 28403 9222
rect 28459 9220 28483 9222
rect 28539 9220 28563 9222
rect 28619 9220 28643 9222
rect 28699 9220 28705 9222
rect 28397 9211 28705 9220
rect 8792 8732 9100 8741
rect 8792 8730 8798 8732
rect 8854 8730 8878 8732
rect 8934 8730 8958 8732
rect 9014 8730 9038 8732
rect 9094 8730 9100 8732
rect 8854 8678 8856 8730
rect 9036 8678 9038 8730
rect 8792 8676 8798 8678
rect 8854 8676 8878 8678
rect 8934 8676 8958 8678
rect 9014 8676 9038 8678
rect 9094 8676 9100 8678
rect 8792 8667 9100 8676
rect 16634 8732 16942 8741
rect 16634 8730 16640 8732
rect 16696 8730 16720 8732
rect 16776 8730 16800 8732
rect 16856 8730 16880 8732
rect 16936 8730 16942 8732
rect 16696 8678 16698 8730
rect 16878 8678 16880 8730
rect 16634 8676 16640 8678
rect 16696 8676 16720 8678
rect 16776 8676 16800 8678
rect 16856 8676 16880 8678
rect 16936 8676 16942 8678
rect 16634 8667 16942 8676
rect 24476 8732 24784 8741
rect 24476 8730 24482 8732
rect 24538 8730 24562 8732
rect 24618 8730 24642 8732
rect 24698 8730 24722 8732
rect 24778 8730 24784 8732
rect 24538 8678 24540 8730
rect 24720 8678 24722 8730
rect 24476 8676 24482 8678
rect 24538 8676 24562 8678
rect 24618 8676 24642 8678
rect 24698 8676 24722 8678
rect 24778 8676 24784 8678
rect 24476 8667 24784 8676
rect 32318 8732 32626 8741
rect 32318 8730 32324 8732
rect 32380 8730 32404 8732
rect 32460 8730 32484 8732
rect 32540 8730 32564 8732
rect 32620 8730 32626 8732
rect 32380 8678 32382 8730
rect 32562 8678 32564 8730
rect 32318 8676 32324 8678
rect 32380 8676 32404 8678
rect 32460 8676 32484 8678
rect 32540 8676 32564 8678
rect 32620 8676 32626 8678
rect 32318 8667 32626 8676
rect 4871 8188 5179 8197
rect 4871 8186 4877 8188
rect 4933 8186 4957 8188
rect 5013 8186 5037 8188
rect 5093 8186 5117 8188
rect 5173 8186 5179 8188
rect 4933 8134 4935 8186
rect 5115 8134 5117 8186
rect 4871 8132 4877 8134
rect 4933 8132 4957 8134
rect 5013 8132 5037 8134
rect 5093 8132 5117 8134
rect 5173 8132 5179 8134
rect 4871 8123 5179 8132
rect 12713 8188 13021 8197
rect 12713 8186 12719 8188
rect 12775 8186 12799 8188
rect 12855 8186 12879 8188
rect 12935 8186 12959 8188
rect 13015 8186 13021 8188
rect 12775 8134 12777 8186
rect 12957 8134 12959 8186
rect 12713 8132 12719 8134
rect 12775 8132 12799 8134
rect 12855 8132 12879 8134
rect 12935 8132 12959 8134
rect 13015 8132 13021 8134
rect 12713 8123 13021 8132
rect 20555 8188 20863 8197
rect 20555 8186 20561 8188
rect 20617 8186 20641 8188
rect 20697 8186 20721 8188
rect 20777 8186 20801 8188
rect 20857 8186 20863 8188
rect 20617 8134 20619 8186
rect 20799 8134 20801 8186
rect 20555 8132 20561 8134
rect 20617 8132 20641 8134
rect 20697 8132 20721 8134
rect 20777 8132 20801 8134
rect 20857 8132 20863 8134
rect 20555 8123 20863 8132
rect 28397 8188 28705 8197
rect 28397 8186 28403 8188
rect 28459 8186 28483 8188
rect 28539 8186 28563 8188
rect 28619 8186 28643 8188
rect 28699 8186 28705 8188
rect 28459 8134 28461 8186
rect 28641 8134 28643 8186
rect 28397 8132 28403 8134
rect 28459 8132 28483 8134
rect 28539 8132 28563 8134
rect 28619 8132 28643 8134
rect 28699 8132 28705 8134
rect 28397 8123 28705 8132
rect 8792 7644 9100 7653
rect 8792 7642 8798 7644
rect 8854 7642 8878 7644
rect 8934 7642 8958 7644
rect 9014 7642 9038 7644
rect 9094 7642 9100 7644
rect 8854 7590 8856 7642
rect 9036 7590 9038 7642
rect 8792 7588 8798 7590
rect 8854 7588 8878 7590
rect 8934 7588 8958 7590
rect 9014 7588 9038 7590
rect 9094 7588 9100 7590
rect 8792 7579 9100 7588
rect 16634 7644 16942 7653
rect 16634 7642 16640 7644
rect 16696 7642 16720 7644
rect 16776 7642 16800 7644
rect 16856 7642 16880 7644
rect 16936 7642 16942 7644
rect 16696 7590 16698 7642
rect 16878 7590 16880 7642
rect 16634 7588 16640 7590
rect 16696 7588 16720 7590
rect 16776 7588 16800 7590
rect 16856 7588 16880 7590
rect 16936 7588 16942 7590
rect 16634 7579 16942 7588
rect 24476 7644 24784 7653
rect 24476 7642 24482 7644
rect 24538 7642 24562 7644
rect 24618 7642 24642 7644
rect 24698 7642 24722 7644
rect 24778 7642 24784 7644
rect 24538 7590 24540 7642
rect 24720 7590 24722 7642
rect 24476 7588 24482 7590
rect 24538 7588 24562 7590
rect 24618 7588 24642 7590
rect 24698 7588 24722 7590
rect 24778 7588 24784 7590
rect 24476 7579 24784 7588
rect 32318 7644 32626 7653
rect 32318 7642 32324 7644
rect 32380 7642 32404 7644
rect 32460 7642 32484 7644
rect 32540 7642 32564 7644
rect 32620 7642 32626 7644
rect 32380 7590 32382 7642
rect 32562 7590 32564 7642
rect 32318 7588 32324 7590
rect 32380 7588 32404 7590
rect 32460 7588 32484 7590
rect 32540 7588 32564 7590
rect 32620 7588 32626 7590
rect 32318 7579 32626 7588
rect 4871 7100 5179 7109
rect 4871 7098 4877 7100
rect 4933 7098 4957 7100
rect 5013 7098 5037 7100
rect 5093 7098 5117 7100
rect 5173 7098 5179 7100
rect 4933 7046 4935 7098
rect 5115 7046 5117 7098
rect 4871 7044 4877 7046
rect 4933 7044 4957 7046
rect 5013 7044 5037 7046
rect 5093 7044 5117 7046
rect 5173 7044 5179 7046
rect 4871 7035 5179 7044
rect 12713 7100 13021 7109
rect 12713 7098 12719 7100
rect 12775 7098 12799 7100
rect 12855 7098 12879 7100
rect 12935 7098 12959 7100
rect 13015 7098 13021 7100
rect 12775 7046 12777 7098
rect 12957 7046 12959 7098
rect 12713 7044 12719 7046
rect 12775 7044 12799 7046
rect 12855 7044 12879 7046
rect 12935 7044 12959 7046
rect 13015 7044 13021 7046
rect 12713 7035 13021 7044
rect 20555 7100 20863 7109
rect 20555 7098 20561 7100
rect 20617 7098 20641 7100
rect 20697 7098 20721 7100
rect 20777 7098 20801 7100
rect 20857 7098 20863 7100
rect 20617 7046 20619 7098
rect 20799 7046 20801 7098
rect 20555 7044 20561 7046
rect 20617 7044 20641 7046
rect 20697 7044 20721 7046
rect 20777 7044 20801 7046
rect 20857 7044 20863 7046
rect 20555 7035 20863 7044
rect 28397 7100 28705 7109
rect 28397 7098 28403 7100
rect 28459 7098 28483 7100
rect 28539 7098 28563 7100
rect 28619 7098 28643 7100
rect 28699 7098 28705 7100
rect 28459 7046 28461 7098
rect 28641 7046 28643 7098
rect 28397 7044 28403 7046
rect 28459 7044 28483 7046
rect 28539 7044 28563 7046
rect 28619 7044 28643 7046
rect 28699 7044 28705 7046
rect 28397 7035 28705 7044
rect 8792 6556 9100 6565
rect 8792 6554 8798 6556
rect 8854 6554 8878 6556
rect 8934 6554 8958 6556
rect 9014 6554 9038 6556
rect 9094 6554 9100 6556
rect 8854 6502 8856 6554
rect 9036 6502 9038 6554
rect 8792 6500 8798 6502
rect 8854 6500 8878 6502
rect 8934 6500 8958 6502
rect 9014 6500 9038 6502
rect 9094 6500 9100 6502
rect 8792 6491 9100 6500
rect 16634 6556 16942 6565
rect 16634 6554 16640 6556
rect 16696 6554 16720 6556
rect 16776 6554 16800 6556
rect 16856 6554 16880 6556
rect 16936 6554 16942 6556
rect 16696 6502 16698 6554
rect 16878 6502 16880 6554
rect 16634 6500 16640 6502
rect 16696 6500 16720 6502
rect 16776 6500 16800 6502
rect 16856 6500 16880 6502
rect 16936 6500 16942 6502
rect 16634 6491 16942 6500
rect 24476 6556 24784 6565
rect 24476 6554 24482 6556
rect 24538 6554 24562 6556
rect 24618 6554 24642 6556
rect 24698 6554 24722 6556
rect 24778 6554 24784 6556
rect 24538 6502 24540 6554
rect 24720 6502 24722 6554
rect 24476 6500 24482 6502
rect 24538 6500 24562 6502
rect 24618 6500 24642 6502
rect 24698 6500 24722 6502
rect 24778 6500 24784 6502
rect 24476 6491 24784 6500
rect 32318 6556 32626 6565
rect 32318 6554 32324 6556
rect 32380 6554 32404 6556
rect 32460 6554 32484 6556
rect 32540 6554 32564 6556
rect 32620 6554 32626 6556
rect 32380 6502 32382 6554
rect 32562 6502 32564 6554
rect 32318 6500 32324 6502
rect 32380 6500 32404 6502
rect 32460 6500 32484 6502
rect 32540 6500 32564 6502
rect 32620 6500 32626 6502
rect 32318 6491 32626 6500
rect 4871 6012 5179 6021
rect 4871 6010 4877 6012
rect 4933 6010 4957 6012
rect 5013 6010 5037 6012
rect 5093 6010 5117 6012
rect 5173 6010 5179 6012
rect 4933 5958 4935 6010
rect 5115 5958 5117 6010
rect 4871 5956 4877 5958
rect 4933 5956 4957 5958
rect 5013 5956 5037 5958
rect 5093 5956 5117 5958
rect 5173 5956 5179 5958
rect 4871 5947 5179 5956
rect 12713 6012 13021 6021
rect 12713 6010 12719 6012
rect 12775 6010 12799 6012
rect 12855 6010 12879 6012
rect 12935 6010 12959 6012
rect 13015 6010 13021 6012
rect 12775 5958 12777 6010
rect 12957 5958 12959 6010
rect 12713 5956 12719 5958
rect 12775 5956 12799 5958
rect 12855 5956 12879 5958
rect 12935 5956 12959 5958
rect 13015 5956 13021 5958
rect 12713 5947 13021 5956
rect 20555 6012 20863 6021
rect 20555 6010 20561 6012
rect 20617 6010 20641 6012
rect 20697 6010 20721 6012
rect 20777 6010 20801 6012
rect 20857 6010 20863 6012
rect 20617 5958 20619 6010
rect 20799 5958 20801 6010
rect 20555 5956 20561 5958
rect 20617 5956 20641 5958
rect 20697 5956 20721 5958
rect 20777 5956 20801 5958
rect 20857 5956 20863 5958
rect 20555 5947 20863 5956
rect 28397 6012 28705 6021
rect 28397 6010 28403 6012
rect 28459 6010 28483 6012
rect 28539 6010 28563 6012
rect 28619 6010 28643 6012
rect 28699 6010 28705 6012
rect 28459 5958 28461 6010
rect 28641 5958 28643 6010
rect 28397 5956 28403 5958
rect 28459 5956 28483 5958
rect 28539 5956 28563 5958
rect 28619 5956 28643 5958
rect 28699 5956 28705 5958
rect 28397 5947 28705 5956
rect 8792 5468 9100 5477
rect 8792 5466 8798 5468
rect 8854 5466 8878 5468
rect 8934 5466 8958 5468
rect 9014 5466 9038 5468
rect 9094 5466 9100 5468
rect 8854 5414 8856 5466
rect 9036 5414 9038 5466
rect 8792 5412 8798 5414
rect 8854 5412 8878 5414
rect 8934 5412 8958 5414
rect 9014 5412 9038 5414
rect 9094 5412 9100 5414
rect 8792 5403 9100 5412
rect 16634 5468 16942 5477
rect 16634 5466 16640 5468
rect 16696 5466 16720 5468
rect 16776 5466 16800 5468
rect 16856 5466 16880 5468
rect 16936 5466 16942 5468
rect 16696 5414 16698 5466
rect 16878 5414 16880 5466
rect 16634 5412 16640 5414
rect 16696 5412 16720 5414
rect 16776 5412 16800 5414
rect 16856 5412 16880 5414
rect 16936 5412 16942 5414
rect 16634 5403 16942 5412
rect 24476 5468 24784 5477
rect 24476 5466 24482 5468
rect 24538 5466 24562 5468
rect 24618 5466 24642 5468
rect 24698 5466 24722 5468
rect 24778 5466 24784 5468
rect 24538 5414 24540 5466
rect 24720 5414 24722 5466
rect 24476 5412 24482 5414
rect 24538 5412 24562 5414
rect 24618 5412 24642 5414
rect 24698 5412 24722 5414
rect 24778 5412 24784 5414
rect 24476 5403 24784 5412
rect 32318 5468 32626 5477
rect 32318 5466 32324 5468
rect 32380 5466 32404 5468
rect 32460 5466 32484 5468
rect 32540 5466 32564 5468
rect 32620 5466 32626 5468
rect 32380 5414 32382 5466
rect 32562 5414 32564 5466
rect 32318 5412 32324 5414
rect 32380 5412 32404 5414
rect 32460 5412 32484 5414
rect 32540 5412 32564 5414
rect 32620 5412 32626 5414
rect 32318 5403 32626 5412
rect 4871 4924 5179 4933
rect 4871 4922 4877 4924
rect 4933 4922 4957 4924
rect 5013 4922 5037 4924
rect 5093 4922 5117 4924
rect 5173 4922 5179 4924
rect 4933 4870 4935 4922
rect 5115 4870 5117 4922
rect 4871 4868 4877 4870
rect 4933 4868 4957 4870
rect 5013 4868 5037 4870
rect 5093 4868 5117 4870
rect 5173 4868 5179 4870
rect 4871 4859 5179 4868
rect 12713 4924 13021 4933
rect 12713 4922 12719 4924
rect 12775 4922 12799 4924
rect 12855 4922 12879 4924
rect 12935 4922 12959 4924
rect 13015 4922 13021 4924
rect 12775 4870 12777 4922
rect 12957 4870 12959 4922
rect 12713 4868 12719 4870
rect 12775 4868 12799 4870
rect 12855 4868 12879 4870
rect 12935 4868 12959 4870
rect 13015 4868 13021 4870
rect 12713 4859 13021 4868
rect 20555 4924 20863 4933
rect 20555 4922 20561 4924
rect 20617 4922 20641 4924
rect 20697 4922 20721 4924
rect 20777 4922 20801 4924
rect 20857 4922 20863 4924
rect 20617 4870 20619 4922
rect 20799 4870 20801 4922
rect 20555 4868 20561 4870
rect 20617 4868 20641 4870
rect 20697 4868 20721 4870
rect 20777 4868 20801 4870
rect 20857 4868 20863 4870
rect 20555 4859 20863 4868
rect 28397 4924 28705 4933
rect 28397 4922 28403 4924
rect 28459 4922 28483 4924
rect 28539 4922 28563 4924
rect 28619 4922 28643 4924
rect 28699 4922 28705 4924
rect 28459 4870 28461 4922
rect 28641 4870 28643 4922
rect 28397 4868 28403 4870
rect 28459 4868 28483 4870
rect 28539 4868 28563 4870
rect 28619 4868 28643 4870
rect 28699 4868 28705 4870
rect 28397 4859 28705 4868
rect 8792 4380 9100 4389
rect 8792 4378 8798 4380
rect 8854 4378 8878 4380
rect 8934 4378 8958 4380
rect 9014 4378 9038 4380
rect 9094 4378 9100 4380
rect 8854 4326 8856 4378
rect 9036 4326 9038 4378
rect 8792 4324 8798 4326
rect 8854 4324 8878 4326
rect 8934 4324 8958 4326
rect 9014 4324 9038 4326
rect 9094 4324 9100 4326
rect 8792 4315 9100 4324
rect 16634 4380 16942 4389
rect 16634 4378 16640 4380
rect 16696 4378 16720 4380
rect 16776 4378 16800 4380
rect 16856 4378 16880 4380
rect 16936 4378 16942 4380
rect 16696 4326 16698 4378
rect 16878 4326 16880 4378
rect 16634 4324 16640 4326
rect 16696 4324 16720 4326
rect 16776 4324 16800 4326
rect 16856 4324 16880 4326
rect 16936 4324 16942 4326
rect 16634 4315 16942 4324
rect 24476 4380 24784 4389
rect 24476 4378 24482 4380
rect 24538 4378 24562 4380
rect 24618 4378 24642 4380
rect 24698 4378 24722 4380
rect 24778 4378 24784 4380
rect 24538 4326 24540 4378
rect 24720 4326 24722 4378
rect 24476 4324 24482 4326
rect 24538 4324 24562 4326
rect 24618 4324 24642 4326
rect 24698 4324 24722 4326
rect 24778 4324 24784 4326
rect 24476 4315 24784 4324
rect 32318 4380 32626 4389
rect 32318 4378 32324 4380
rect 32380 4378 32404 4380
rect 32460 4378 32484 4380
rect 32540 4378 32564 4380
rect 32620 4378 32626 4380
rect 32380 4326 32382 4378
rect 32562 4326 32564 4378
rect 32318 4324 32324 4326
rect 32380 4324 32404 4326
rect 32460 4324 32484 4326
rect 32540 4324 32564 4326
rect 32620 4324 32626 4326
rect 32318 4315 32626 4324
rect 4871 3836 5179 3845
rect 4871 3834 4877 3836
rect 4933 3834 4957 3836
rect 5013 3834 5037 3836
rect 5093 3834 5117 3836
rect 5173 3834 5179 3836
rect 4933 3782 4935 3834
rect 5115 3782 5117 3834
rect 4871 3780 4877 3782
rect 4933 3780 4957 3782
rect 5013 3780 5037 3782
rect 5093 3780 5117 3782
rect 5173 3780 5179 3782
rect 4871 3771 5179 3780
rect 12713 3836 13021 3845
rect 12713 3834 12719 3836
rect 12775 3834 12799 3836
rect 12855 3834 12879 3836
rect 12935 3834 12959 3836
rect 13015 3834 13021 3836
rect 12775 3782 12777 3834
rect 12957 3782 12959 3834
rect 12713 3780 12719 3782
rect 12775 3780 12799 3782
rect 12855 3780 12879 3782
rect 12935 3780 12959 3782
rect 13015 3780 13021 3782
rect 12713 3771 13021 3780
rect 20555 3836 20863 3845
rect 20555 3834 20561 3836
rect 20617 3834 20641 3836
rect 20697 3834 20721 3836
rect 20777 3834 20801 3836
rect 20857 3834 20863 3836
rect 20617 3782 20619 3834
rect 20799 3782 20801 3834
rect 20555 3780 20561 3782
rect 20617 3780 20641 3782
rect 20697 3780 20721 3782
rect 20777 3780 20801 3782
rect 20857 3780 20863 3782
rect 20555 3771 20863 3780
rect 28397 3836 28705 3845
rect 28397 3834 28403 3836
rect 28459 3834 28483 3836
rect 28539 3834 28563 3836
rect 28619 3834 28643 3836
rect 28699 3834 28705 3836
rect 28459 3782 28461 3834
rect 28641 3782 28643 3834
rect 28397 3780 28403 3782
rect 28459 3780 28483 3782
rect 28539 3780 28563 3782
rect 28619 3780 28643 3782
rect 28699 3780 28705 3782
rect 28397 3771 28705 3780
rect 8792 3292 9100 3301
rect 8792 3290 8798 3292
rect 8854 3290 8878 3292
rect 8934 3290 8958 3292
rect 9014 3290 9038 3292
rect 9094 3290 9100 3292
rect 8854 3238 8856 3290
rect 9036 3238 9038 3290
rect 8792 3236 8798 3238
rect 8854 3236 8878 3238
rect 8934 3236 8958 3238
rect 9014 3236 9038 3238
rect 9094 3236 9100 3238
rect 8792 3227 9100 3236
rect 16634 3292 16942 3301
rect 16634 3290 16640 3292
rect 16696 3290 16720 3292
rect 16776 3290 16800 3292
rect 16856 3290 16880 3292
rect 16936 3290 16942 3292
rect 16696 3238 16698 3290
rect 16878 3238 16880 3290
rect 16634 3236 16640 3238
rect 16696 3236 16720 3238
rect 16776 3236 16800 3238
rect 16856 3236 16880 3238
rect 16936 3236 16942 3238
rect 16634 3227 16942 3236
rect 24476 3292 24784 3301
rect 24476 3290 24482 3292
rect 24538 3290 24562 3292
rect 24618 3290 24642 3292
rect 24698 3290 24722 3292
rect 24778 3290 24784 3292
rect 24538 3238 24540 3290
rect 24720 3238 24722 3290
rect 24476 3236 24482 3238
rect 24538 3236 24562 3238
rect 24618 3236 24642 3238
rect 24698 3236 24722 3238
rect 24778 3236 24784 3238
rect 24476 3227 24784 3236
rect 32318 3292 32626 3301
rect 32318 3290 32324 3292
rect 32380 3290 32404 3292
rect 32460 3290 32484 3292
rect 32540 3290 32564 3292
rect 32620 3290 32626 3292
rect 32380 3238 32382 3290
rect 32562 3238 32564 3290
rect 32318 3236 32324 3238
rect 32380 3236 32404 3238
rect 32460 3236 32484 3238
rect 32540 3236 32564 3238
rect 32620 3236 32626 3238
rect 32318 3227 32626 3236
rect 4871 2748 5179 2757
rect 4871 2746 4877 2748
rect 4933 2746 4957 2748
rect 5013 2746 5037 2748
rect 5093 2746 5117 2748
rect 5173 2746 5179 2748
rect 4933 2694 4935 2746
rect 5115 2694 5117 2746
rect 4871 2692 4877 2694
rect 4933 2692 4957 2694
rect 5013 2692 5037 2694
rect 5093 2692 5117 2694
rect 5173 2692 5179 2694
rect 4871 2683 5179 2692
rect 12713 2748 13021 2757
rect 12713 2746 12719 2748
rect 12775 2746 12799 2748
rect 12855 2746 12879 2748
rect 12935 2746 12959 2748
rect 13015 2746 13021 2748
rect 12775 2694 12777 2746
rect 12957 2694 12959 2746
rect 12713 2692 12719 2694
rect 12775 2692 12799 2694
rect 12855 2692 12879 2694
rect 12935 2692 12959 2694
rect 13015 2692 13021 2694
rect 12713 2683 13021 2692
rect 20555 2748 20863 2757
rect 20555 2746 20561 2748
rect 20617 2746 20641 2748
rect 20697 2746 20721 2748
rect 20777 2746 20801 2748
rect 20857 2746 20863 2748
rect 20617 2694 20619 2746
rect 20799 2694 20801 2746
rect 20555 2692 20561 2694
rect 20617 2692 20641 2694
rect 20697 2692 20721 2694
rect 20777 2692 20801 2694
rect 20857 2692 20863 2694
rect 20555 2683 20863 2692
rect 28397 2748 28705 2757
rect 28397 2746 28403 2748
rect 28459 2746 28483 2748
rect 28539 2746 28563 2748
rect 28619 2746 28643 2748
rect 28699 2746 28705 2748
rect 28459 2694 28461 2746
rect 28641 2694 28643 2746
rect 28397 2692 28403 2694
rect 28459 2692 28483 2694
rect 28539 2692 28563 2694
rect 28619 2692 28643 2694
rect 28699 2692 28705 2694
rect 28397 2683 28705 2692
rect 8792 2204 9100 2213
rect 8792 2202 8798 2204
rect 8854 2202 8878 2204
rect 8934 2202 8958 2204
rect 9014 2202 9038 2204
rect 9094 2202 9100 2204
rect 8854 2150 8856 2202
rect 9036 2150 9038 2202
rect 8792 2148 8798 2150
rect 8854 2148 8878 2150
rect 8934 2148 8958 2150
rect 9014 2148 9038 2150
rect 9094 2148 9100 2150
rect 8792 2139 9100 2148
rect 16634 2204 16942 2213
rect 16634 2202 16640 2204
rect 16696 2202 16720 2204
rect 16776 2202 16800 2204
rect 16856 2202 16880 2204
rect 16936 2202 16942 2204
rect 16696 2150 16698 2202
rect 16878 2150 16880 2202
rect 16634 2148 16640 2150
rect 16696 2148 16720 2150
rect 16776 2148 16800 2150
rect 16856 2148 16880 2150
rect 16936 2148 16942 2150
rect 16634 2139 16942 2148
rect 24476 2204 24784 2213
rect 24476 2202 24482 2204
rect 24538 2202 24562 2204
rect 24618 2202 24642 2204
rect 24698 2202 24722 2204
rect 24778 2202 24784 2204
rect 24538 2150 24540 2202
rect 24720 2150 24722 2202
rect 24476 2148 24482 2150
rect 24538 2148 24562 2150
rect 24618 2148 24642 2150
rect 24698 2148 24722 2150
rect 24778 2148 24784 2150
rect 24476 2139 24784 2148
rect 32318 2204 32626 2213
rect 32318 2202 32324 2204
rect 32380 2202 32404 2204
rect 32460 2202 32484 2204
rect 32540 2202 32564 2204
rect 32620 2202 32626 2204
rect 32380 2150 32382 2202
rect 32562 2150 32564 2202
rect 32318 2148 32324 2150
rect 32380 2148 32404 2150
rect 32460 2148 32484 2150
rect 32540 2148 32564 2150
rect 32620 2148 32626 2150
rect 32318 2139 32626 2148
rect 4871 1660 5179 1669
rect 4871 1658 4877 1660
rect 4933 1658 4957 1660
rect 5013 1658 5037 1660
rect 5093 1658 5117 1660
rect 5173 1658 5179 1660
rect 4933 1606 4935 1658
rect 5115 1606 5117 1658
rect 4871 1604 4877 1606
rect 4933 1604 4957 1606
rect 5013 1604 5037 1606
rect 5093 1604 5117 1606
rect 5173 1604 5179 1606
rect 4871 1595 5179 1604
rect 12713 1660 13021 1669
rect 12713 1658 12719 1660
rect 12775 1658 12799 1660
rect 12855 1658 12879 1660
rect 12935 1658 12959 1660
rect 13015 1658 13021 1660
rect 12775 1606 12777 1658
rect 12957 1606 12959 1658
rect 12713 1604 12719 1606
rect 12775 1604 12799 1606
rect 12855 1604 12879 1606
rect 12935 1604 12959 1606
rect 13015 1604 13021 1606
rect 12713 1595 13021 1604
rect 20555 1660 20863 1669
rect 20555 1658 20561 1660
rect 20617 1658 20641 1660
rect 20697 1658 20721 1660
rect 20777 1658 20801 1660
rect 20857 1658 20863 1660
rect 20617 1606 20619 1658
rect 20799 1606 20801 1658
rect 20555 1604 20561 1606
rect 20617 1604 20641 1606
rect 20697 1604 20721 1606
rect 20777 1604 20801 1606
rect 20857 1604 20863 1606
rect 20555 1595 20863 1604
rect 28397 1660 28705 1669
rect 28397 1658 28403 1660
rect 28459 1658 28483 1660
rect 28539 1658 28563 1660
rect 28619 1658 28643 1660
rect 28699 1658 28705 1660
rect 28459 1606 28461 1658
rect 28641 1606 28643 1658
rect 28397 1604 28403 1606
rect 28459 1604 28483 1606
rect 28539 1604 28563 1606
rect 28619 1604 28643 1606
rect 28699 1604 28705 1606
rect 28397 1595 28705 1604
rect 8792 1116 9100 1125
rect 8792 1114 8798 1116
rect 8854 1114 8878 1116
rect 8934 1114 8958 1116
rect 9014 1114 9038 1116
rect 9094 1114 9100 1116
rect 8854 1062 8856 1114
rect 9036 1062 9038 1114
rect 8792 1060 8798 1062
rect 8854 1060 8878 1062
rect 8934 1060 8958 1062
rect 9014 1060 9038 1062
rect 9094 1060 9100 1062
rect 8792 1051 9100 1060
rect 16634 1116 16942 1125
rect 16634 1114 16640 1116
rect 16696 1114 16720 1116
rect 16776 1114 16800 1116
rect 16856 1114 16880 1116
rect 16936 1114 16942 1116
rect 16696 1062 16698 1114
rect 16878 1062 16880 1114
rect 16634 1060 16640 1062
rect 16696 1060 16720 1062
rect 16776 1060 16800 1062
rect 16856 1060 16880 1062
rect 16936 1060 16942 1062
rect 16634 1051 16942 1060
rect 24476 1116 24784 1125
rect 24476 1114 24482 1116
rect 24538 1114 24562 1116
rect 24618 1114 24642 1116
rect 24698 1114 24722 1116
rect 24778 1114 24784 1116
rect 24538 1062 24540 1114
rect 24720 1062 24722 1114
rect 24476 1060 24482 1062
rect 24538 1060 24562 1062
rect 24618 1060 24642 1062
rect 24698 1060 24722 1062
rect 24778 1060 24784 1062
rect 24476 1051 24784 1060
rect 32318 1116 32626 1125
rect 32318 1114 32324 1116
rect 32380 1114 32404 1116
rect 32460 1114 32484 1116
rect 32540 1114 32564 1116
rect 32620 1114 32626 1116
rect 32380 1062 32382 1114
rect 32562 1062 32564 1114
rect 32318 1060 32324 1062
rect 32380 1060 32404 1062
rect 32460 1060 32484 1062
rect 32540 1060 32564 1062
rect 32620 1060 32626 1062
rect 32318 1051 32626 1060
<< via2 >>
rect 9126 21392 9182 21448
rect 9678 21392 9734 21448
rect 11058 21392 11114 21448
rect 11886 21392 11942 21448
rect 12806 21392 12862 21448
rect 14002 21392 14058 21448
rect 15566 21392 15622 21448
rect 15750 21392 15806 21448
rect 17498 21392 17554 21448
rect 19246 21392 19302 21448
rect 19522 21392 19578 21448
rect 21730 21392 21786 21448
rect 22926 21392 22982 21448
rect 23662 21392 23718 21448
rect 24398 21392 24454 21448
rect 25870 21392 25926 21448
rect 27434 21392 27490 21448
rect 28814 21392 28870 21448
rect 30286 21392 30342 21448
rect 5170 20848 5226 20904
rect 2134 20460 2190 20496
rect 2134 20440 2136 20460
rect 2136 20440 2188 20460
rect 2188 20440 2190 20460
rect 2778 20460 2834 20496
rect 2778 20440 2780 20460
rect 2780 20440 2832 20460
rect 2832 20440 2834 20460
rect 3422 20460 3478 20496
rect 3422 20440 3424 20460
rect 3424 20440 3476 20460
rect 3476 20440 3478 20460
rect 4526 20460 4582 20496
rect 8798 20698 8854 20700
rect 8878 20698 8934 20700
rect 8958 20698 9014 20700
rect 9038 20698 9094 20700
rect 8798 20646 8844 20698
rect 8844 20646 8854 20698
rect 8878 20646 8908 20698
rect 8908 20646 8920 20698
rect 8920 20646 8934 20698
rect 8958 20646 8972 20698
rect 8972 20646 8984 20698
rect 8984 20646 9014 20698
rect 9038 20646 9048 20698
rect 9048 20646 9094 20698
rect 8798 20644 8854 20646
rect 8878 20644 8934 20646
rect 8958 20644 9014 20646
rect 9038 20644 9094 20646
rect 4526 20440 4528 20460
rect 4528 20440 4580 20460
rect 4580 20440 4582 20460
rect 5998 20460 6054 20496
rect 5998 20440 6000 20460
rect 6000 20440 6052 20460
rect 6052 20440 6054 20460
rect 4877 20154 4933 20156
rect 4957 20154 5013 20156
rect 5037 20154 5093 20156
rect 5117 20154 5173 20156
rect 4877 20102 4923 20154
rect 4923 20102 4933 20154
rect 4957 20102 4987 20154
rect 4987 20102 4999 20154
rect 4999 20102 5013 20154
rect 5037 20102 5051 20154
rect 5051 20102 5063 20154
rect 5063 20102 5093 20154
rect 5117 20102 5127 20154
rect 5127 20102 5173 20154
rect 4877 20100 4933 20102
rect 4957 20100 5013 20102
rect 5037 20100 5093 20102
rect 5117 20100 5173 20102
rect 1582 20052 1638 20088
rect 1582 20032 1584 20052
rect 1584 20032 1636 20052
rect 1636 20032 1638 20052
rect 6734 20052 6790 20088
rect 6734 20032 6736 20052
rect 6736 20032 6788 20052
rect 6788 20032 6790 20052
rect 7470 20052 7526 20088
rect 7470 20032 7472 20052
rect 7472 20032 7524 20052
rect 7524 20032 7526 20052
rect 8206 20052 8262 20088
rect 8206 20032 8208 20052
rect 8208 20032 8260 20052
rect 8260 20032 8262 20052
rect 8798 19610 8854 19612
rect 8878 19610 8934 19612
rect 8958 19610 9014 19612
rect 9038 19610 9094 19612
rect 8798 19558 8844 19610
rect 8844 19558 8854 19610
rect 8878 19558 8908 19610
rect 8908 19558 8920 19610
rect 8920 19558 8934 19610
rect 8958 19558 8972 19610
rect 8972 19558 8984 19610
rect 8984 19558 9014 19610
rect 9038 19558 9048 19610
rect 9048 19558 9094 19610
rect 8798 19556 8854 19558
rect 8878 19556 8934 19558
rect 8958 19556 9014 19558
rect 9038 19556 9094 19558
rect 10138 20052 10194 20088
rect 10138 20032 10140 20052
rect 10140 20032 10192 20052
rect 10192 20032 10194 20052
rect 4877 19066 4933 19068
rect 4957 19066 5013 19068
rect 5037 19066 5093 19068
rect 5117 19066 5173 19068
rect 4877 19014 4923 19066
rect 4923 19014 4933 19066
rect 4957 19014 4987 19066
rect 4987 19014 4999 19066
rect 4999 19014 5013 19066
rect 5037 19014 5051 19066
rect 5051 19014 5063 19066
rect 5063 19014 5093 19066
rect 5117 19014 5127 19066
rect 5127 19014 5173 19066
rect 4877 19012 4933 19014
rect 4957 19012 5013 19014
rect 5037 19012 5093 19014
rect 5117 19012 5173 19014
rect 8798 18522 8854 18524
rect 8878 18522 8934 18524
rect 8958 18522 9014 18524
rect 9038 18522 9094 18524
rect 8798 18470 8844 18522
rect 8844 18470 8854 18522
rect 8878 18470 8908 18522
rect 8908 18470 8920 18522
rect 8920 18470 8934 18522
rect 8958 18470 8972 18522
rect 8972 18470 8984 18522
rect 8984 18470 9014 18522
rect 9038 18470 9048 18522
rect 9048 18470 9094 18522
rect 8798 18468 8854 18470
rect 8878 18468 8934 18470
rect 8958 18468 9014 18470
rect 9038 18468 9094 18470
rect 4877 17978 4933 17980
rect 4957 17978 5013 17980
rect 5037 17978 5093 17980
rect 5117 17978 5173 17980
rect 4877 17926 4923 17978
rect 4923 17926 4933 17978
rect 4957 17926 4987 17978
rect 4987 17926 4999 17978
rect 4999 17926 5013 17978
rect 5037 17926 5051 17978
rect 5051 17926 5063 17978
rect 5063 17926 5093 17978
rect 5117 17926 5127 17978
rect 5127 17926 5173 17978
rect 4877 17924 4933 17926
rect 4957 17924 5013 17926
rect 5037 17924 5093 17926
rect 5117 17924 5173 17926
rect 8798 17434 8854 17436
rect 8878 17434 8934 17436
rect 8958 17434 9014 17436
rect 9038 17434 9094 17436
rect 8798 17382 8844 17434
rect 8844 17382 8854 17434
rect 8878 17382 8908 17434
rect 8908 17382 8920 17434
rect 8920 17382 8934 17434
rect 8958 17382 8972 17434
rect 8972 17382 8984 17434
rect 8984 17382 9014 17434
rect 9038 17382 9048 17434
rect 9048 17382 9094 17434
rect 8798 17380 8854 17382
rect 8878 17380 8934 17382
rect 8958 17380 9014 17382
rect 9038 17380 9094 17382
rect 4877 16890 4933 16892
rect 4957 16890 5013 16892
rect 5037 16890 5093 16892
rect 5117 16890 5173 16892
rect 4877 16838 4923 16890
rect 4923 16838 4933 16890
rect 4957 16838 4987 16890
rect 4987 16838 4999 16890
rect 4999 16838 5013 16890
rect 5037 16838 5051 16890
rect 5051 16838 5063 16890
rect 5063 16838 5093 16890
rect 5117 16838 5127 16890
rect 5127 16838 5173 16890
rect 4877 16836 4933 16838
rect 4957 16836 5013 16838
rect 5037 16836 5093 16838
rect 5117 16836 5173 16838
rect 8798 16346 8854 16348
rect 8878 16346 8934 16348
rect 8958 16346 9014 16348
rect 9038 16346 9094 16348
rect 8798 16294 8844 16346
rect 8844 16294 8854 16346
rect 8878 16294 8908 16346
rect 8908 16294 8920 16346
rect 8920 16294 8934 16346
rect 8958 16294 8972 16346
rect 8972 16294 8984 16346
rect 8984 16294 9014 16346
rect 9038 16294 9048 16346
rect 9048 16294 9094 16346
rect 8798 16292 8854 16294
rect 8878 16292 8934 16294
rect 8958 16292 9014 16294
rect 9038 16292 9094 16294
rect 4877 15802 4933 15804
rect 4957 15802 5013 15804
rect 5037 15802 5093 15804
rect 5117 15802 5173 15804
rect 4877 15750 4923 15802
rect 4923 15750 4933 15802
rect 4957 15750 4987 15802
rect 4987 15750 4999 15802
rect 4999 15750 5013 15802
rect 5037 15750 5051 15802
rect 5051 15750 5063 15802
rect 5063 15750 5093 15802
rect 5117 15750 5127 15802
rect 5127 15750 5173 15802
rect 4877 15748 4933 15750
rect 4957 15748 5013 15750
rect 5037 15748 5093 15750
rect 5117 15748 5173 15750
rect 8798 15258 8854 15260
rect 8878 15258 8934 15260
rect 8958 15258 9014 15260
rect 9038 15258 9094 15260
rect 8798 15206 8844 15258
rect 8844 15206 8854 15258
rect 8878 15206 8908 15258
rect 8908 15206 8920 15258
rect 8920 15206 8934 15258
rect 8958 15206 8972 15258
rect 8972 15206 8984 15258
rect 8984 15206 9014 15258
rect 9038 15206 9048 15258
rect 9048 15206 9094 15258
rect 8798 15204 8854 15206
rect 8878 15204 8934 15206
rect 8958 15204 9014 15206
rect 9038 15204 9094 15206
rect 4877 14714 4933 14716
rect 4957 14714 5013 14716
rect 5037 14714 5093 14716
rect 5117 14714 5173 14716
rect 4877 14662 4923 14714
rect 4923 14662 4933 14714
rect 4957 14662 4987 14714
rect 4987 14662 4999 14714
rect 4999 14662 5013 14714
rect 5037 14662 5051 14714
rect 5051 14662 5063 14714
rect 5063 14662 5093 14714
rect 5117 14662 5127 14714
rect 5127 14662 5173 14714
rect 4877 14660 4933 14662
rect 4957 14660 5013 14662
rect 5037 14660 5093 14662
rect 5117 14660 5173 14662
rect 8798 14170 8854 14172
rect 8878 14170 8934 14172
rect 8958 14170 9014 14172
rect 9038 14170 9094 14172
rect 8798 14118 8844 14170
rect 8844 14118 8854 14170
rect 8878 14118 8908 14170
rect 8908 14118 8920 14170
rect 8920 14118 8934 14170
rect 8958 14118 8972 14170
rect 8972 14118 8984 14170
rect 8984 14118 9014 14170
rect 9038 14118 9048 14170
rect 9048 14118 9094 14170
rect 8798 14116 8854 14118
rect 8878 14116 8934 14118
rect 8958 14116 9014 14118
rect 9038 14116 9094 14118
rect 4877 13626 4933 13628
rect 4957 13626 5013 13628
rect 5037 13626 5093 13628
rect 5117 13626 5173 13628
rect 4877 13574 4923 13626
rect 4923 13574 4933 13626
rect 4957 13574 4987 13626
rect 4987 13574 4999 13626
rect 4999 13574 5013 13626
rect 5037 13574 5051 13626
rect 5051 13574 5063 13626
rect 5063 13574 5093 13626
rect 5117 13574 5127 13626
rect 5127 13574 5173 13626
rect 4877 13572 4933 13574
rect 4957 13572 5013 13574
rect 5037 13572 5093 13574
rect 5117 13572 5173 13574
rect 8798 13082 8854 13084
rect 8878 13082 8934 13084
rect 8958 13082 9014 13084
rect 9038 13082 9094 13084
rect 8798 13030 8844 13082
rect 8844 13030 8854 13082
rect 8878 13030 8908 13082
rect 8908 13030 8920 13082
rect 8920 13030 8934 13082
rect 8958 13030 8972 13082
rect 8972 13030 8984 13082
rect 8984 13030 9014 13082
rect 9038 13030 9048 13082
rect 9048 13030 9094 13082
rect 8798 13028 8854 13030
rect 8878 13028 8934 13030
rect 8958 13028 9014 13030
rect 9038 13028 9094 13030
rect 12622 20304 12678 20360
rect 13818 21256 13874 21312
rect 12719 20154 12775 20156
rect 12799 20154 12855 20156
rect 12879 20154 12935 20156
rect 12959 20154 13015 20156
rect 12719 20102 12765 20154
rect 12765 20102 12775 20154
rect 12799 20102 12829 20154
rect 12829 20102 12841 20154
rect 12841 20102 12855 20154
rect 12879 20102 12893 20154
rect 12893 20102 12905 20154
rect 12905 20102 12935 20154
rect 12959 20102 12969 20154
rect 12969 20102 13015 20154
rect 12719 20100 12775 20102
rect 12799 20100 12855 20102
rect 12879 20100 12935 20102
rect 12959 20100 13015 20102
rect 12719 19066 12775 19068
rect 12799 19066 12855 19068
rect 12879 19066 12935 19068
rect 12959 19066 13015 19068
rect 12719 19014 12765 19066
rect 12765 19014 12775 19066
rect 12799 19014 12829 19066
rect 12829 19014 12841 19066
rect 12841 19014 12855 19066
rect 12879 19014 12893 19066
rect 12893 19014 12905 19066
rect 12905 19014 12935 19066
rect 12959 19014 12969 19066
rect 12969 19014 13015 19066
rect 12719 19012 12775 19014
rect 12799 19012 12855 19014
rect 12879 19012 12935 19014
rect 12959 19012 13015 19014
rect 16640 20698 16696 20700
rect 16720 20698 16776 20700
rect 16800 20698 16856 20700
rect 16880 20698 16936 20700
rect 16640 20646 16686 20698
rect 16686 20646 16696 20698
rect 16720 20646 16750 20698
rect 16750 20646 16762 20698
rect 16762 20646 16776 20698
rect 16800 20646 16814 20698
rect 16814 20646 16826 20698
rect 16826 20646 16856 20698
rect 16880 20646 16890 20698
rect 16890 20646 16936 20698
rect 16640 20644 16696 20646
rect 16720 20644 16776 20646
rect 16800 20644 16856 20646
rect 16880 20644 16936 20646
rect 16640 19610 16696 19612
rect 16720 19610 16776 19612
rect 16800 19610 16856 19612
rect 16880 19610 16936 19612
rect 16640 19558 16686 19610
rect 16686 19558 16696 19610
rect 16720 19558 16750 19610
rect 16750 19558 16762 19610
rect 16762 19558 16776 19610
rect 16800 19558 16814 19610
rect 16814 19558 16826 19610
rect 16826 19558 16856 19610
rect 16880 19558 16890 19610
rect 16890 19558 16936 19610
rect 16640 19556 16696 19558
rect 16720 19556 16776 19558
rect 16800 19556 16856 19558
rect 16880 19556 16936 19558
rect 17866 21256 17922 21312
rect 16640 18522 16696 18524
rect 16720 18522 16776 18524
rect 16800 18522 16856 18524
rect 16880 18522 16936 18524
rect 16640 18470 16686 18522
rect 16686 18470 16696 18522
rect 16720 18470 16750 18522
rect 16750 18470 16762 18522
rect 16762 18470 16776 18522
rect 16800 18470 16814 18522
rect 16814 18470 16826 18522
rect 16826 18470 16856 18522
rect 16880 18470 16890 18522
rect 16890 18470 16936 18522
rect 16640 18468 16696 18470
rect 16720 18468 16776 18470
rect 16800 18468 16856 18470
rect 16880 18468 16936 18470
rect 12719 17978 12775 17980
rect 12799 17978 12855 17980
rect 12879 17978 12935 17980
rect 12959 17978 13015 17980
rect 12719 17926 12765 17978
rect 12765 17926 12775 17978
rect 12799 17926 12829 17978
rect 12829 17926 12841 17978
rect 12841 17926 12855 17978
rect 12879 17926 12893 17978
rect 12893 17926 12905 17978
rect 12905 17926 12935 17978
rect 12959 17926 12969 17978
rect 12969 17926 13015 17978
rect 12719 17924 12775 17926
rect 12799 17924 12855 17926
rect 12879 17924 12935 17926
rect 12959 17924 13015 17926
rect 16640 17434 16696 17436
rect 16720 17434 16776 17436
rect 16800 17434 16856 17436
rect 16880 17434 16936 17436
rect 16640 17382 16686 17434
rect 16686 17382 16696 17434
rect 16720 17382 16750 17434
rect 16750 17382 16762 17434
rect 16762 17382 16776 17434
rect 16800 17382 16814 17434
rect 16814 17382 16826 17434
rect 16826 17382 16856 17434
rect 16880 17382 16890 17434
rect 16890 17382 16936 17434
rect 16640 17380 16696 17382
rect 16720 17380 16776 17382
rect 16800 17380 16856 17382
rect 16880 17380 16936 17382
rect 12719 16890 12775 16892
rect 12799 16890 12855 16892
rect 12879 16890 12935 16892
rect 12959 16890 13015 16892
rect 12719 16838 12765 16890
rect 12765 16838 12775 16890
rect 12799 16838 12829 16890
rect 12829 16838 12841 16890
rect 12841 16838 12855 16890
rect 12879 16838 12893 16890
rect 12893 16838 12905 16890
rect 12905 16838 12935 16890
rect 12959 16838 12969 16890
rect 12969 16838 13015 16890
rect 12719 16836 12775 16838
rect 12799 16836 12855 16838
rect 12879 16836 12935 16838
rect 12959 16836 13015 16838
rect 16640 16346 16696 16348
rect 16720 16346 16776 16348
rect 16800 16346 16856 16348
rect 16880 16346 16936 16348
rect 16640 16294 16686 16346
rect 16686 16294 16696 16346
rect 16720 16294 16750 16346
rect 16750 16294 16762 16346
rect 16762 16294 16776 16346
rect 16800 16294 16814 16346
rect 16814 16294 16826 16346
rect 16826 16294 16856 16346
rect 16880 16294 16890 16346
rect 16890 16294 16936 16346
rect 16640 16292 16696 16294
rect 16720 16292 16776 16294
rect 16800 16292 16856 16294
rect 16880 16292 16936 16294
rect 21226 21216 21296 21276
rect 20902 20848 20958 20904
rect 20561 20154 20617 20156
rect 20641 20154 20697 20156
rect 20721 20154 20777 20156
rect 20801 20154 20857 20156
rect 20561 20102 20607 20154
rect 20607 20102 20617 20154
rect 20641 20102 20671 20154
rect 20671 20102 20683 20154
rect 20683 20102 20697 20154
rect 20721 20102 20735 20154
rect 20735 20102 20747 20154
rect 20747 20102 20777 20154
rect 20801 20102 20811 20154
rect 20811 20102 20857 20154
rect 20561 20100 20617 20102
rect 20641 20100 20697 20102
rect 20721 20100 20777 20102
rect 20801 20100 20857 20102
rect 20810 19932 20812 19952
rect 20812 19932 20864 19952
rect 20864 19932 20866 19952
rect 20810 19896 20866 19932
rect 12719 15802 12775 15804
rect 12799 15802 12855 15804
rect 12879 15802 12935 15804
rect 12959 15802 13015 15804
rect 12719 15750 12765 15802
rect 12765 15750 12775 15802
rect 12799 15750 12829 15802
rect 12829 15750 12841 15802
rect 12841 15750 12855 15802
rect 12879 15750 12893 15802
rect 12893 15750 12905 15802
rect 12905 15750 12935 15802
rect 12959 15750 12969 15802
rect 12969 15750 13015 15802
rect 12719 15748 12775 15750
rect 12799 15748 12855 15750
rect 12879 15748 12935 15750
rect 12959 15748 13015 15750
rect 16640 15258 16696 15260
rect 16720 15258 16776 15260
rect 16800 15258 16856 15260
rect 16880 15258 16936 15260
rect 16640 15206 16686 15258
rect 16686 15206 16696 15258
rect 16720 15206 16750 15258
rect 16750 15206 16762 15258
rect 16762 15206 16776 15258
rect 16800 15206 16814 15258
rect 16814 15206 16826 15258
rect 16826 15206 16856 15258
rect 16880 15206 16890 15258
rect 16890 15206 16936 15258
rect 16640 15204 16696 15206
rect 16720 15204 16776 15206
rect 16800 15204 16856 15206
rect 16880 15204 16936 15206
rect 12719 14714 12775 14716
rect 12799 14714 12855 14716
rect 12879 14714 12935 14716
rect 12959 14714 13015 14716
rect 12719 14662 12765 14714
rect 12765 14662 12775 14714
rect 12799 14662 12829 14714
rect 12829 14662 12841 14714
rect 12841 14662 12855 14714
rect 12879 14662 12893 14714
rect 12893 14662 12905 14714
rect 12905 14662 12935 14714
rect 12959 14662 12969 14714
rect 12969 14662 13015 14714
rect 12719 14660 12775 14662
rect 12799 14660 12855 14662
rect 12879 14660 12935 14662
rect 12959 14660 13015 14662
rect 20626 19252 20628 19272
rect 20628 19252 20680 19272
rect 20680 19252 20682 19272
rect 20626 19216 20682 19252
rect 20561 19066 20617 19068
rect 20641 19066 20697 19068
rect 20721 19066 20777 19068
rect 20801 19066 20857 19068
rect 20561 19014 20607 19066
rect 20607 19014 20617 19066
rect 20641 19014 20671 19066
rect 20671 19014 20683 19066
rect 20683 19014 20697 19066
rect 20721 19014 20735 19066
rect 20735 19014 20747 19066
rect 20747 19014 20777 19066
rect 20801 19014 20811 19066
rect 20811 19014 20857 19066
rect 20561 19012 20617 19014
rect 20641 19012 20697 19014
rect 20721 19012 20777 19014
rect 20801 19012 20857 19014
rect 20561 17978 20617 17980
rect 20641 17978 20697 17980
rect 20721 17978 20777 17980
rect 20801 17978 20857 17980
rect 20561 17926 20607 17978
rect 20607 17926 20617 17978
rect 20641 17926 20671 17978
rect 20671 17926 20683 17978
rect 20683 17926 20697 17978
rect 20721 17926 20735 17978
rect 20735 17926 20747 17978
rect 20747 17926 20777 17978
rect 20801 17926 20811 17978
rect 20811 17926 20857 17978
rect 20561 17924 20617 17926
rect 20641 17924 20697 17926
rect 20721 17924 20777 17926
rect 20801 17924 20857 17926
rect 20561 16890 20617 16892
rect 20641 16890 20697 16892
rect 20721 16890 20777 16892
rect 20801 16890 20857 16892
rect 20561 16838 20607 16890
rect 20607 16838 20617 16890
rect 20641 16838 20671 16890
rect 20671 16838 20683 16890
rect 20683 16838 20697 16890
rect 20721 16838 20735 16890
rect 20735 16838 20747 16890
rect 20747 16838 20777 16890
rect 20801 16838 20811 16890
rect 20811 16838 20857 16890
rect 20561 16836 20617 16838
rect 20641 16836 20697 16838
rect 20721 16836 20777 16838
rect 20801 16836 20857 16838
rect 21178 19896 21234 19952
rect 20561 15802 20617 15804
rect 20641 15802 20697 15804
rect 20721 15802 20777 15804
rect 20801 15802 20857 15804
rect 20561 15750 20607 15802
rect 20607 15750 20617 15802
rect 20641 15750 20671 15802
rect 20671 15750 20683 15802
rect 20683 15750 20697 15802
rect 20721 15750 20735 15802
rect 20735 15750 20747 15802
rect 20747 15750 20777 15802
rect 20801 15750 20811 15802
rect 20811 15750 20857 15802
rect 20561 15748 20617 15750
rect 20641 15748 20697 15750
rect 20721 15748 20777 15750
rect 20801 15748 20857 15750
rect 20561 14714 20617 14716
rect 20641 14714 20697 14716
rect 20721 14714 20777 14716
rect 20801 14714 20857 14716
rect 20561 14662 20607 14714
rect 20607 14662 20617 14714
rect 20641 14662 20671 14714
rect 20671 14662 20683 14714
rect 20683 14662 20697 14714
rect 20721 14662 20735 14714
rect 20735 14662 20747 14714
rect 20747 14662 20777 14714
rect 20801 14662 20811 14714
rect 20811 14662 20857 14714
rect 20561 14660 20617 14662
rect 20641 14660 20697 14662
rect 20721 14660 20777 14662
rect 20801 14660 20857 14662
rect 16640 14170 16696 14172
rect 16720 14170 16776 14172
rect 16800 14170 16856 14172
rect 16880 14170 16936 14172
rect 16640 14118 16686 14170
rect 16686 14118 16696 14170
rect 16720 14118 16750 14170
rect 16750 14118 16762 14170
rect 16762 14118 16776 14170
rect 16800 14118 16814 14170
rect 16814 14118 16826 14170
rect 16826 14118 16856 14170
rect 16880 14118 16890 14170
rect 16890 14118 16936 14170
rect 16640 14116 16696 14118
rect 16720 14116 16776 14118
rect 16800 14116 16856 14118
rect 16880 14116 16936 14118
rect 12719 13626 12775 13628
rect 12799 13626 12855 13628
rect 12879 13626 12935 13628
rect 12959 13626 13015 13628
rect 12719 13574 12765 13626
rect 12765 13574 12775 13626
rect 12799 13574 12829 13626
rect 12829 13574 12841 13626
rect 12841 13574 12855 13626
rect 12879 13574 12893 13626
rect 12893 13574 12905 13626
rect 12905 13574 12935 13626
rect 12959 13574 12969 13626
rect 12969 13574 13015 13626
rect 12719 13572 12775 13574
rect 12799 13572 12855 13574
rect 12879 13572 12935 13574
rect 12959 13572 13015 13574
rect 16640 13082 16696 13084
rect 16720 13082 16776 13084
rect 16800 13082 16856 13084
rect 16880 13082 16936 13084
rect 16640 13030 16686 13082
rect 16686 13030 16696 13082
rect 16720 13030 16750 13082
rect 16750 13030 16762 13082
rect 16762 13030 16776 13082
rect 16800 13030 16814 13082
rect 16814 13030 16826 13082
rect 16826 13030 16856 13082
rect 16880 13030 16890 13082
rect 16890 13030 16936 13082
rect 16640 13028 16696 13030
rect 16720 13028 16776 13030
rect 16800 13028 16856 13030
rect 16880 13028 16936 13030
rect 4877 12538 4933 12540
rect 4957 12538 5013 12540
rect 5037 12538 5093 12540
rect 5117 12538 5173 12540
rect 4877 12486 4923 12538
rect 4923 12486 4933 12538
rect 4957 12486 4987 12538
rect 4987 12486 4999 12538
rect 4999 12486 5013 12538
rect 5037 12486 5051 12538
rect 5051 12486 5063 12538
rect 5063 12486 5093 12538
rect 5117 12486 5127 12538
rect 5127 12486 5173 12538
rect 4877 12484 4933 12486
rect 4957 12484 5013 12486
rect 5037 12484 5093 12486
rect 5117 12484 5173 12486
rect 12719 12538 12775 12540
rect 12799 12538 12855 12540
rect 12879 12538 12935 12540
rect 12959 12538 13015 12540
rect 12719 12486 12765 12538
rect 12765 12486 12775 12538
rect 12799 12486 12829 12538
rect 12829 12486 12841 12538
rect 12841 12486 12855 12538
rect 12879 12486 12893 12538
rect 12893 12486 12905 12538
rect 12905 12486 12935 12538
rect 12959 12486 12969 12538
rect 12969 12486 13015 12538
rect 12719 12484 12775 12486
rect 12799 12484 12855 12486
rect 12879 12484 12935 12486
rect 12959 12484 13015 12486
rect 20561 13626 20617 13628
rect 20641 13626 20697 13628
rect 20721 13626 20777 13628
rect 20801 13626 20857 13628
rect 20561 13574 20607 13626
rect 20607 13574 20617 13626
rect 20641 13574 20671 13626
rect 20671 13574 20683 13626
rect 20683 13574 20697 13626
rect 20721 13574 20735 13626
rect 20735 13574 20747 13626
rect 20747 13574 20777 13626
rect 20801 13574 20811 13626
rect 20811 13574 20857 13626
rect 20561 13572 20617 13574
rect 20641 13572 20697 13574
rect 20721 13572 20777 13574
rect 20801 13572 20857 13574
rect 20561 12538 20617 12540
rect 20641 12538 20697 12540
rect 20721 12538 20777 12540
rect 20801 12538 20857 12540
rect 20561 12486 20607 12538
rect 20607 12486 20617 12538
rect 20641 12486 20671 12538
rect 20671 12486 20683 12538
rect 20683 12486 20697 12538
rect 20721 12486 20735 12538
rect 20735 12486 20747 12538
rect 20747 12486 20777 12538
rect 20801 12486 20811 12538
rect 20811 12486 20857 12538
rect 20561 12484 20617 12486
rect 20641 12484 20697 12486
rect 20721 12484 20777 12486
rect 20801 12484 20857 12486
rect 21822 19488 21878 19544
rect 22006 19216 22062 19272
rect 23570 19488 23626 19544
rect 24482 20698 24538 20700
rect 24562 20698 24618 20700
rect 24642 20698 24698 20700
rect 24722 20698 24778 20700
rect 24482 20646 24528 20698
rect 24528 20646 24538 20698
rect 24562 20646 24592 20698
rect 24592 20646 24604 20698
rect 24604 20646 24618 20698
rect 24642 20646 24656 20698
rect 24656 20646 24668 20698
rect 24668 20646 24698 20698
rect 24722 20646 24732 20698
rect 24732 20646 24778 20698
rect 24482 20644 24538 20646
rect 24562 20644 24618 20646
rect 24642 20644 24698 20646
rect 24722 20644 24778 20646
rect 24766 20440 24822 20496
rect 27342 20984 27398 21040
rect 28630 20984 28686 21040
rect 24482 19610 24538 19612
rect 24562 19610 24618 19612
rect 24642 19610 24698 19612
rect 24722 19610 24778 19612
rect 24482 19558 24528 19610
rect 24528 19558 24538 19610
rect 24562 19558 24592 19610
rect 24592 19558 24604 19610
rect 24604 19558 24618 19610
rect 24642 19558 24656 19610
rect 24656 19558 24668 19610
rect 24668 19558 24698 19610
rect 24722 19558 24732 19610
rect 24732 19558 24778 19610
rect 24482 19556 24538 19558
rect 24562 19556 24618 19558
rect 24642 19556 24698 19558
rect 24722 19556 24778 19558
rect 24482 18522 24538 18524
rect 24562 18522 24618 18524
rect 24642 18522 24698 18524
rect 24722 18522 24778 18524
rect 24482 18470 24528 18522
rect 24528 18470 24538 18522
rect 24562 18470 24592 18522
rect 24592 18470 24604 18522
rect 24604 18470 24618 18522
rect 24642 18470 24656 18522
rect 24656 18470 24668 18522
rect 24668 18470 24698 18522
rect 24722 18470 24732 18522
rect 24732 18470 24778 18522
rect 24482 18468 24538 18470
rect 24562 18468 24618 18470
rect 24642 18468 24698 18470
rect 24722 18468 24778 18470
rect 24482 17434 24538 17436
rect 24562 17434 24618 17436
rect 24642 17434 24698 17436
rect 24722 17434 24778 17436
rect 24482 17382 24528 17434
rect 24528 17382 24538 17434
rect 24562 17382 24592 17434
rect 24592 17382 24604 17434
rect 24604 17382 24618 17434
rect 24642 17382 24656 17434
rect 24656 17382 24668 17434
rect 24668 17382 24698 17434
rect 24722 17382 24732 17434
rect 24732 17382 24778 17434
rect 24482 17380 24538 17382
rect 24562 17380 24618 17382
rect 24642 17380 24698 17382
rect 24722 17380 24778 17382
rect 24482 16346 24538 16348
rect 24562 16346 24618 16348
rect 24642 16346 24698 16348
rect 24722 16346 24778 16348
rect 24482 16294 24528 16346
rect 24528 16294 24538 16346
rect 24562 16294 24592 16346
rect 24592 16294 24604 16346
rect 24604 16294 24618 16346
rect 24642 16294 24656 16346
rect 24656 16294 24668 16346
rect 24668 16294 24698 16346
rect 24722 16294 24732 16346
rect 24732 16294 24778 16346
rect 24482 16292 24538 16294
rect 24562 16292 24618 16294
rect 24642 16292 24698 16294
rect 24722 16292 24778 16294
rect 24482 15258 24538 15260
rect 24562 15258 24618 15260
rect 24642 15258 24698 15260
rect 24722 15258 24778 15260
rect 24482 15206 24528 15258
rect 24528 15206 24538 15258
rect 24562 15206 24592 15258
rect 24592 15206 24604 15258
rect 24604 15206 24618 15258
rect 24642 15206 24656 15258
rect 24656 15206 24668 15258
rect 24668 15206 24698 15258
rect 24722 15206 24732 15258
rect 24732 15206 24778 15258
rect 24482 15204 24538 15206
rect 24562 15204 24618 15206
rect 24642 15204 24698 15206
rect 24722 15204 24778 15206
rect 24482 14170 24538 14172
rect 24562 14170 24618 14172
rect 24642 14170 24698 14172
rect 24722 14170 24778 14172
rect 24482 14118 24528 14170
rect 24528 14118 24538 14170
rect 24562 14118 24592 14170
rect 24592 14118 24604 14170
rect 24604 14118 24618 14170
rect 24642 14118 24656 14170
rect 24656 14118 24668 14170
rect 24668 14118 24698 14170
rect 24722 14118 24732 14170
rect 24732 14118 24778 14170
rect 24482 14116 24538 14118
rect 24562 14116 24618 14118
rect 24642 14116 24698 14118
rect 24722 14116 24778 14118
rect 28403 20154 28459 20156
rect 28483 20154 28539 20156
rect 28563 20154 28619 20156
rect 28643 20154 28699 20156
rect 28403 20102 28449 20154
rect 28449 20102 28459 20154
rect 28483 20102 28513 20154
rect 28513 20102 28525 20154
rect 28525 20102 28539 20154
rect 28563 20102 28577 20154
rect 28577 20102 28589 20154
rect 28589 20102 28619 20154
rect 28643 20102 28653 20154
rect 28653 20102 28699 20154
rect 28403 20100 28459 20102
rect 28483 20100 28539 20102
rect 28563 20100 28619 20102
rect 28643 20100 28699 20102
rect 29918 20984 29974 21040
rect 33614 21208 33696 21280
rect 32324 20698 32380 20700
rect 32404 20698 32460 20700
rect 32484 20698 32540 20700
rect 32564 20698 32620 20700
rect 32324 20646 32370 20698
rect 32370 20646 32380 20698
rect 32404 20646 32434 20698
rect 32434 20646 32446 20698
rect 32446 20646 32460 20698
rect 32484 20646 32498 20698
rect 32498 20646 32510 20698
rect 32510 20646 32540 20698
rect 32564 20646 32574 20698
rect 32574 20646 32620 20698
rect 32324 20644 32380 20646
rect 32404 20644 32460 20646
rect 32484 20644 32540 20646
rect 32564 20644 32620 20646
rect 28403 19066 28459 19068
rect 28483 19066 28539 19068
rect 28563 19066 28619 19068
rect 28643 19066 28699 19068
rect 28403 19014 28449 19066
rect 28449 19014 28459 19066
rect 28483 19014 28513 19066
rect 28513 19014 28525 19066
rect 28525 19014 28539 19066
rect 28563 19014 28577 19066
rect 28577 19014 28589 19066
rect 28589 19014 28619 19066
rect 28643 19014 28653 19066
rect 28653 19014 28699 19066
rect 28403 19012 28459 19014
rect 28483 19012 28539 19014
rect 28563 19012 28619 19014
rect 28643 19012 28699 19014
rect 28403 17978 28459 17980
rect 28483 17978 28539 17980
rect 28563 17978 28619 17980
rect 28643 17978 28699 17980
rect 28403 17926 28449 17978
rect 28449 17926 28459 17978
rect 28483 17926 28513 17978
rect 28513 17926 28525 17978
rect 28525 17926 28539 17978
rect 28563 17926 28577 17978
rect 28577 17926 28589 17978
rect 28589 17926 28619 17978
rect 28643 17926 28653 17978
rect 28653 17926 28699 17978
rect 28403 17924 28459 17926
rect 28483 17924 28539 17926
rect 28563 17924 28619 17926
rect 28643 17924 28699 17926
rect 28403 16890 28459 16892
rect 28483 16890 28539 16892
rect 28563 16890 28619 16892
rect 28643 16890 28699 16892
rect 28403 16838 28449 16890
rect 28449 16838 28459 16890
rect 28483 16838 28513 16890
rect 28513 16838 28525 16890
rect 28525 16838 28539 16890
rect 28563 16838 28577 16890
rect 28577 16838 28589 16890
rect 28589 16838 28619 16890
rect 28643 16838 28653 16890
rect 28653 16838 28699 16890
rect 28403 16836 28459 16838
rect 28483 16836 28539 16838
rect 28563 16836 28619 16838
rect 28643 16836 28699 16838
rect 28403 15802 28459 15804
rect 28483 15802 28539 15804
rect 28563 15802 28619 15804
rect 28643 15802 28699 15804
rect 28403 15750 28449 15802
rect 28449 15750 28459 15802
rect 28483 15750 28513 15802
rect 28513 15750 28525 15802
rect 28525 15750 28539 15802
rect 28563 15750 28577 15802
rect 28577 15750 28589 15802
rect 28589 15750 28619 15802
rect 28643 15750 28653 15802
rect 28653 15750 28699 15802
rect 28403 15748 28459 15750
rect 28483 15748 28539 15750
rect 28563 15748 28619 15750
rect 28643 15748 28699 15750
rect 28403 14714 28459 14716
rect 28483 14714 28539 14716
rect 28563 14714 28619 14716
rect 28643 14714 28699 14716
rect 28403 14662 28449 14714
rect 28449 14662 28459 14714
rect 28483 14662 28513 14714
rect 28513 14662 28525 14714
rect 28525 14662 28539 14714
rect 28563 14662 28577 14714
rect 28577 14662 28589 14714
rect 28589 14662 28619 14714
rect 28643 14662 28653 14714
rect 28653 14662 28699 14714
rect 28403 14660 28459 14662
rect 28483 14660 28539 14662
rect 28563 14660 28619 14662
rect 28643 14660 28699 14662
rect 32324 19610 32380 19612
rect 32404 19610 32460 19612
rect 32484 19610 32540 19612
rect 32564 19610 32620 19612
rect 32324 19558 32370 19610
rect 32370 19558 32380 19610
rect 32404 19558 32434 19610
rect 32434 19558 32446 19610
rect 32446 19558 32460 19610
rect 32484 19558 32498 19610
rect 32498 19558 32510 19610
rect 32510 19558 32540 19610
rect 32564 19558 32574 19610
rect 32574 19558 32620 19610
rect 32324 19556 32380 19558
rect 32404 19556 32460 19558
rect 32484 19556 32540 19558
rect 32564 19556 32620 19558
rect 32324 18522 32380 18524
rect 32404 18522 32460 18524
rect 32484 18522 32540 18524
rect 32564 18522 32620 18524
rect 32324 18470 32370 18522
rect 32370 18470 32380 18522
rect 32404 18470 32434 18522
rect 32434 18470 32446 18522
rect 32446 18470 32460 18522
rect 32484 18470 32498 18522
rect 32498 18470 32510 18522
rect 32510 18470 32540 18522
rect 32564 18470 32574 18522
rect 32574 18470 32620 18522
rect 32324 18468 32380 18470
rect 32404 18468 32460 18470
rect 32484 18468 32540 18470
rect 32564 18468 32620 18470
rect 32324 17434 32380 17436
rect 32404 17434 32460 17436
rect 32484 17434 32540 17436
rect 32564 17434 32620 17436
rect 32324 17382 32370 17434
rect 32370 17382 32380 17434
rect 32404 17382 32434 17434
rect 32434 17382 32446 17434
rect 32446 17382 32460 17434
rect 32484 17382 32498 17434
rect 32498 17382 32510 17434
rect 32510 17382 32540 17434
rect 32564 17382 32574 17434
rect 32574 17382 32620 17434
rect 32324 17380 32380 17382
rect 32404 17380 32460 17382
rect 32484 17380 32540 17382
rect 32564 17380 32620 17382
rect 32324 16346 32380 16348
rect 32404 16346 32460 16348
rect 32484 16346 32540 16348
rect 32564 16346 32620 16348
rect 32324 16294 32370 16346
rect 32370 16294 32380 16346
rect 32404 16294 32434 16346
rect 32434 16294 32446 16346
rect 32446 16294 32460 16346
rect 32484 16294 32498 16346
rect 32498 16294 32510 16346
rect 32510 16294 32540 16346
rect 32564 16294 32574 16346
rect 32574 16294 32620 16346
rect 32324 16292 32380 16294
rect 32404 16292 32460 16294
rect 32484 16292 32540 16294
rect 32564 16292 32620 16294
rect 32324 15258 32380 15260
rect 32404 15258 32460 15260
rect 32484 15258 32540 15260
rect 32564 15258 32620 15260
rect 32324 15206 32370 15258
rect 32370 15206 32380 15258
rect 32404 15206 32434 15258
rect 32434 15206 32446 15258
rect 32446 15206 32460 15258
rect 32484 15206 32498 15258
rect 32498 15206 32510 15258
rect 32510 15206 32540 15258
rect 32564 15206 32574 15258
rect 32574 15206 32620 15258
rect 32324 15204 32380 15206
rect 32404 15204 32460 15206
rect 32484 15204 32540 15206
rect 32564 15204 32620 15206
rect 32324 14170 32380 14172
rect 32404 14170 32460 14172
rect 32484 14170 32540 14172
rect 32564 14170 32620 14172
rect 32324 14118 32370 14170
rect 32370 14118 32380 14170
rect 32404 14118 32434 14170
rect 32434 14118 32446 14170
rect 32446 14118 32460 14170
rect 32484 14118 32498 14170
rect 32498 14118 32510 14170
rect 32510 14118 32540 14170
rect 32564 14118 32574 14170
rect 32574 14118 32620 14170
rect 32324 14116 32380 14118
rect 32404 14116 32460 14118
rect 32484 14116 32540 14118
rect 32564 14116 32620 14118
rect 28403 13626 28459 13628
rect 28483 13626 28539 13628
rect 28563 13626 28619 13628
rect 28643 13626 28699 13628
rect 28403 13574 28449 13626
rect 28449 13574 28459 13626
rect 28483 13574 28513 13626
rect 28513 13574 28525 13626
rect 28525 13574 28539 13626
rect 28563 13574 28577 13626
rect 28577 13574 28589 13626
rect 28589 13574 28619 13626
rect 28643 13574 28653 13626
rect 28653 13574 28699 13626
rect 28403 13572 28459 13574
rect 28483 13572 28539 13574
rect 28563 13572 28619 13574
rect 28643 13572 28699 13574
rect 24482 13082 24538 13084
rect 24562 13082 24618 13084
rect 24642 13082 24698 13084
rect 24722 13082 24778 13084
rect 24482 13030 24528 13082
rect 24528 13030 24538 13082
rect 24562 13030 24592 13082
rect 24592 13030 24604 13082
rect 24604 13030 24618 13082
rect 24642 13030 24656 13082
rect 24656 13030 24668 13082
rect 24668 13030 24698 13082
rect 24722 13030 24732 13082
rect 24732 13030 24778 13082
rect 24482 13028 24538 13030
rect 24562 13028 24618 13030
rect 24642 13028 24698 13030
rect 24722 13028 24778 13030
rect 32324 13082 32380 13084
rect 32404 13082 32460 13084
rect 32484 13082 32540 13084
rect 32564 13082 32620 13084
rect 32324 13030 32370 13082
rect 32370 13030 32380 13082
rect 32404 13030 32434 13082
rect 32434 13030 32446 13082
rect 32446 13030 32460 13082
rect 32484 13030 32498 13082
rect 32498 13030 32510 13082
rect 32510 13030 32540 13082
rect 32564 13030 32574 13082
rect 32574 13030 32620 13082
rect 32324 13028 32380 13030
rect 32404 13028 32460 13030
rect 32484 13028 32540 13030
rect 32564 13028 32620 13030
rect 28403 12538 28459 12540
rect 28483 12538 28539 12540
rect 28563 12538 28619 12540
rect 28643 12538 28699 12540
rect 28403 12486 28449 12538
rect 28449 12486 28459 12538
rect 28483 12486 28513 12538
rect 28513 12486 28525 12538
rect 28525 12486 28539 12538
rect 28563 12486 28577 12538
rect 28577 12486 28589 12538
rect 28589 12486 28619 12538
rect 28643 12486 28653 12538
rect 28653 12486 28699 12538
rect 28403 12484 28459 12486
rect 28483 12484 28539 12486
rect 28563 12484 28619 12486
rect 28643 12484 28699 12486
rect 8798 11994 8854 11996
rect 8878 11994 8934 11996
rect 8958 11994 9014 11996
rect 9038 11994 9094 11996
rect 8798 11942 8844 11994
rect 8844 11942 8854 11994
rect 8878 11942 8908 11994
rect 8908 11942 8920 11994
rect 8920 11942 8934 11994
rect 8958 11942 8972 11994
rect 8972 11942 8984 11994
rect 8984 11942 9014 11994
rect 9038 11942 9048 11994
rect 9048 11942 9094 11994
rect 8798 11940 8854 11942
rect 8878 11940 8934 11942
rect 8958 11940 9014 11942
rect 9038 11940 9094 11942
rect 16640 11994 16696 11996
rect 16720 11994 16776 11996
rect 16800 11994 16856 11996
rect 16880 11994 16936 11996
rect 16640 11942 16686 11994
rect 16686 11942 16696 11994
rect 16720 11942 16750 11994
rect 16750 11942 16762 11994
rect 16762 11942 16776 11994
rect 16800 11942 16814 11994
rect 16814 11942 16826 11994
rect 16826 11942 16856 11994
rect 16880 11942 16890 11994
rect 16890 11942 16936 11994
rect 16640 11940 16696 11942
rect 16720 11940 16776 11942
rect 16800 11940 16856 11942
rect 16880 11940 16936 11942
rect 24482 11994 24538 11996
rect 24562 11994 24618 11996
rect 24642 11994 24698 11996
rect 24722 11994 24778 11996
rect 24482 11942 24528 11994
rect 24528 11942 24538 11994
rect 24562 11942 24592 11994
rect 24592 11942 24604 11994
rect 24604 11942 24618 11994
rect 24642 11942 24656 11994
rect 24656 11942 24668 11994
rect 24668 11942 24698 11994
rect 24722 11942 24732 11994
rect 24732 11942 24778 11994
rect 24482 11940 24538 11942
rect 24562 11940 24618 11942
rect 24642 11940 24698 11942
rect 24722 11940 24778 11942
rect 32324 11994 32380 11996
rect 32404 11994 32460 11996
rect 32484 11994 32540 11996
rect 32564 11994 32620 11996
rect 32324 11942 32370 11994
rect 32370 11942 32380 11994
rect 32404 11942 32434 11994
rect 32434 11942 32446 11994
rect 32446 11942 32460 11994
rect 32484 11942 32498 11994
rect 32498 11942 32510 11994
rect 32510 11942 32540 11994
rect 32564 11942 32574 11994
rect 32574 11942 32620 11994
rect 32324 11940 32380 11942
rect 32404 11940 32460 11942
rect 32484 11940 32540 11942
rect 32564 11940 32620 11942
rect 4877 11450 4933 11452
rect 4957 11450 5013 11452
rect 5037 11450 5093 11452
rect 5117 11450 5173 11452
rect 4877 11398 4923 11450
rect 4923 11398 4933 11450
rect 4957 11398 4987 11450
rect 4987 11398 4999 11450
rect 4999 11398 5013 11450
rect 5037 11398 5051 11450
rect 5051 11398 5063 11450
rect 5063 11398 5093 11450
rect 5117 11398 5127 11450
rect 5127 11398 5173 11450
rect 4877 11396 4933 11398
rect 4957 11396 5013 11398
rect 5037 11396 5093 11398
rect 5117 11396 5173 11398
rect 12719 11450 12775 11452
rect 12799 11450 12855 11452
rect 12879 11450 12935 11452
rect 12959 11450 13015 11452
rect 12719 11398 12765 11450
rect 12765 11398 12775 11450
rect 12799 11398 12829 11450
rect 12829 11398 12841 11450
rect 12841 11398 12855 11450
rect 12879 11398 12893 11450
rect 12893 11398 12905 11450
rect 12905 11398 12935 11450
rect 12959 11398 12969 11450
rect 12969 11398 13015 11450
rect 12719 11396 12775 11398
rect 12799 11396 12855 11398
rect 12879 11396 12935 11398
rect 12959 11396 13015 11398
rect 20561 11450 20617 11452
rect 20641 11450 20697 11452
rect 20721 11450 20777 11452
rect 20801 11450 20857 11452
rect 20561 11398 20607 11450
rect 20607 11398 20617 11450
rect 20641 11398 20671 11450
rect 20671 11398 20683 11450
rect 20683 11398 20697 11450
rect 20721 11398 20735 11450
rect 20735 11398 20747 11450
rect 20747 11398 20777 11450
rect 20801 11398 20811 11450
rect 20811 11398 20857 11450
rect 20561 11396 20617 11398
rect 20641 11396 20697 11398
rect 20721 11396 20777 11398
rect 20801 11396 20857 11398
rect 28403 11450 28459 11452
rect 28483 11450 28539 11452
rect 28563 11450 28619 11452
rect 28643 11450 28699 11452
rect 28403 11398 28449 11450
rect 28449 11398 28459 11450
rect 28483 11398 28513 11450
rect 28513 11398 28525 11450
rect 28525 11398 28539 11450
rect 28563 11398 28577 11450
rect 28577 11398 28589 11450
rect 28589 11398 28619 11450
rect 28643 11398 28653 11450
rect 28653 11398 28699 11450
rect 28403 11396 28459 11398
rect 28483 11396 28539 11398
rect 28563 11396 28619 11398
rect 28643 11396 28699 11398
rect 8798 10906 8854 10908
rect 8878 10906 8934 10908
rect 8958 10906 9014 10908
rect 9038 10906 9094 10908
rect 8798 10854 8844 10906
rect 8844 10854 8854 10906
rect 8878 10854 8908 10906
rect 8908 10854 8920 10906
rect 8920 10854 8934 10906
rect 8958 10854 8972 10906
rect 8972 10854 8984 10906
rect 8984 10854 9014 10906
rect 9038 10854 9048 10906
rect 9048 10854 9094 10906
rect 8798 10852 8854 10854
rect 8878 10852 8934 10854
rect 8958 10852 9014 10854
rect 9038 10852 9094 10854
rect 16640 10906 16696 10908
rect 16720 10906 16776 10908
rect 16800 10906 16856 10908
rect 16880 10906 16936 10908
rect 16640 10854 16686 10906
rect 16686 10854 16696 10906
rect 16720 10854 16750 10906
rect 16750 10854 16762 10906
rect 16762 10854 16776 10906
rect 16800 10854 16814 10906
rect 16814 10854 16826 10906
rect 16826 10854 16856 10906
rect 16880 10854 16890 10906
rect 16890 10854 16936 10906
rect 16640 10852 16696 10854
rect 16720 10852 16776 10854
rect 16800 10852 16856 10854
rect 16880 10852 16936 10854
rect 24482 10906 24538 10908
rect 24562 10906 24618 10908
rect 24642 10906 24698 10908
rect 24722 10906 24778 10908
rect 24482 10854 24528 10906
rect 24528 10854 24538 10906
rect 24562 10854 24592 10906
rect 24592 10854 24604 10906
rect 24604 10854 24618 10906
rect 24642 10854 24656 10906
rect 24656 10854 24668 10906
rect 24668 10854 24698 10906
rect 24722 10854 24732 10906
rect 24732 10854 24778 10906
rect 24482 10852 24538 10854
rect 24562 10852 24618 10854
rect 24642 10852 24698 10854
rect 24722 10852 24778 10854
rect 32324 10906 32380 10908
rect 32404 10906 32460 10908
rect 32484 10906 32540 10908
rect 32564 10906 32620 10908
rect 32324 10854 32370 10906
rect 32370 10854 32380 10906
rect 32404 10854 32434 10906
rect 32434 10854 32446 10906
rect 32446 10854 32460 10906
rect 32484 10854 32498 10906
rect 32498 10854 32510 10906
rect 32510 10854 32540 10906
rect 32564 10854 32574 10906
rect 32574 10854 32620 10906
rect 32324 10852 32380 10854
rect 32404 10852 32460 10854
rect 32484 10852 32540 10854
rect 32564 10852 32620 10854
rect 4877 10362 4933 10364
rect 4957 10362 5013 10364
rect 5037 10362 5093 10364
rect 5117 10362 5173 10364
rect 4877 10310 4923 10362
rect 4923 10310 4933 10362
rect 4957 10310 4987 10362
rect 4987 10310 4999 10362
rect 4999 10310 5013 10362
rect 5037 10310 5051 10362
rect 5051 10310 5063 10362
rect 5063 10310 5093 10362
rect 5117 10310 5127 10362
rect 5127 10310 5173 10362
rect 4877 10308 4933 10310
rect 4957 10308 5013 10310
rect 5037 10308 5093 10310
rect 5117 10308 5173 10310
rect 12719 10362 12775 10364
rect 12799 10362 12855 10364
rect 12879 10362 12935 10364
rect 12959 10362 13015 10364
rect 12719 10310 12765 10362
rect 12765 10310 12775 10362
rect 12799 10310 12829 10362
rect 12829 10310 12841 10362
rect 12841 10310 12855 10362
rect 12879 10310 12893 10362
rect 12893 10310 12905 10362
rect 12905 10310 12935 10362
rect 12959 10310 12969 10362
rect 12969 10310 13015 10362
rect 12719 10308 12775 10310
rect 12799 10308 12855 10310
rect 12879 10308 12935 10310
rect 12959 10308 13015 10310
rect 20561 10362 20617 10364
rect 20641 10362 20697 10364
rect 20721 10362 20777 10364
rect 20801 10362 20857 10364
rect 20561 10310 20607 10362
rect 20607 10310 20617 10362
rect 20641 10310 20671 10362
rect 20671 10310 20683 10362
rect 20683 10310 20697 10362
rect 20721 10310 20735 10362
rect 20735 10310 20747 10362
rect 20747 10310 20777 10362
rect 20801 10310 20811 10362
rect 20811 10310 20857 10362
rect 20561 10308 20617 10310
rect 20641 10308 20697 10310
rect 20721 10308 20777 10310
rect 20801 10308 20857 10310
rect 28403 10362 28459 10364
rect 28483 10362 28539 10364
rect 28563 10362 28619 10364
rect 28643 10362 28699 10364
rect 28403 10310 28449 10362
rect 28449 10310 28459 10362
rect 28483 10310 28513 10362
rect 28513 10310 28525 10362
rect 28525 10310 28539 10362
rect 28563 10310 28577 10362
rect 28577 10310 28589 10362
rect 28589 10310 28619 10362
rect 28643 10310 28653 10362
rect 28653 10310 28699 10362
rect 28403 10308 28459 10310
rect 28483 10308 28539 10310
rect 28563 10308 28619 10310
rect 28643 10308 28699 10310
rect 8798 9818 8854 9820
rect 8878 9818 8934 9820
rect 8958 9818 9014 9820
rect 9038 9818 9094 9820
rect 8798 9766 8844 9818
rect 8844 9766 8854 9818
rect 8878 9766 8908 9818
rect 8908 9766 8920 9818
rect 8920 9766 8934 9818
rect 8958 9766 8972 9818
rect 8972 9766 8984 9818
rect 8984 9766 9014 9818
rect 9038 9766 9048 9818
rect 9048 9766 9094 9818
rect 8798 9764 8854 9766
rect 8878 9764 8934 9766
rect 8958 9764 9014 9766
rect 9038 9764 9094 9766
rect 16640 9818 16696 9820
rect 16720 9818 16776 9820
rect 16800 9818 16856 9820
rect 16880 9818 16936 9820
rect 16640 9766 16686 9818
rect 16686 9766 16696 9818
rect 16720 9766 16750 9818
rect 16750 9766 16762 9818
rect 16762 9766 16776 9818
rect 16800 9766 16814 9818
rect 16814 9766 16826 9818
rect 16826 9766 16856 9818
rect 16880 9766 16890 9818
rect 16890 9766 16936 9818
rect 16640 9764 16696 9766
rect 16720 9764 16776 9766
rect 16800 9764 16856 9766
rect 16880 9764 16936 9766
rect 24482 9818 24538 9820
rect 24562 9818 24618 9820
rect 24642 9818 24698 9820
rect 24722 9818 24778 9820
rect 24482 9766 24528 9818
rect 24528 9766 24538 9818
rect 24562 9766 24592 9818
rect 24592 9766 24604 9818
rect 24604 9766 24618 9818
rect 24642 9766 24656 9818
rect 24656 9766 24668 9818
rect 24668 9766 24698 9818
rect 24722 9766 24732 9818
rect 24732 9766 24778 9818
rect 24482 9764 24538 9766
rect 24562 9764 24618 9766
rect 24642 9764 24698 9766
rect 24722 9764 24778 9766
rect 32324 9818 32380 9820
rect 32404 9818 32460 9820
rect 32484 9818 32540 9820
rect 32564 9818 32620 9820
rect 32324 9766 32370 9818
rect 32370 9766 32380 9818
rect 32404 9766 32434 9818
rect 32434 9766 32446 9818
rect 32446 9766 32460 9818
rect 32484 9766 32498 9818
rect 32498 9766 32510 9818
rect 32510 9766 32540 9818
rect 32564 9766 32574 9818
rect 32574 9766 32620 9818
rect 32324 9764 32380 9766
rect 32404 9764 32460 9766
rect 32484 9764 32540 9766
rect 32564 9764 32620 9766
rect 4877 9274 4933 9276
rect 4957 9274 5013 9276
rect 5037 9274 5093 9276
rect 5117 9274 5173 9276
rect 4877 9222 4923 9274
rect 4923 9222 4933 9274
rect 4957 9222 4987 9274
rect 4987 9222 4999 9274
rect 4999 9222 5013 9274
rect 5037 9222 5051 9274
rect 5051 9222 5063 9274
rect 5063 9222 5093 9274
rect 5117 9222 5127 9274
rect 5127 9222 5173 9274
rect 4877 9220 4933 9222
rect 4957 9220 5013 9222
rect 5037 9220 5093 9222
rect 5117 9220 5173 9222
rect 12719 9274 12775 9276
rect 12799 9274 12855 9276
rect 12879 9274 12935 9276
rect 12959 9274 13015 9276
rect 12719 9222 12765 9274
rect 12765 9222 12775 9274
rect 12799 9222 12829 9274
rect 12829 9222 12841 9274
rect 12841 9222 12855 9274
rect 12879 9222 12893 9274
rect 12893 9222 12905 9274
rect 12905 9222 12935 9274
rect 12959 9222 12969 9274
rect 12969 9222 13015 9274
rect 12719 9220 12775 9222
rect 12799 9220 12855 9222
rect 12879 9220 12935 9222
rect 12959 9220 13015 9222
rect 20561 9274 20617 9276
rect 20641 9274 20697 9276
rect 20721 9274 20777 9276
rect 20801 9274 20857 9276
rect 20561 9222 20607 9274
rect 20607 9222 20617 9274
rect 20641 9222 20671 9274
rect 20671 9222 20683 9274
rect 20683 9222 20697 9274
rect 20721 9222 20735 9274
rect 20735 9222 20747 9274
rect 20747 9222 20777 9274
rect 20801 9222 20811 9274
rect 20811 9222 20857 9274
rect 20561 9220 20617 9222
rect 20641 9220 20697 9222
rect 20721 9220 20777 9222
rect 20801 9220 20857 9222
rect 28403 9274 28459 9276
rect 28483 9274 28539 9276
rect 28563 9274 28619 9276
rect 28643 9274 28699 9276
rect 28403 9222 28449 9274
rect 28449 9222 28459 9274
rect 28483 9222 28513 9274
rect 28513 9222 28525 9274
rect 28525 9222 28539 9274
rect 28563 9222 28577 9274
rect 28577 9222 28589 9274
rect 28589 9222 28619 9274
rect 28643 9222 28653 9274
rect 28653 9222 28699 9274
rect 28403 9220 28459 9222
rect 28483 9220 28539 9222
rect 28563 9220 28619 9222
rect 28643 9220 28699 9222
rect 8798 8730 8854 8732
rect 8878 8730 8934 8732
rect 8958 8730 9014 8732
rect 9038 8730 9094 8732
rect 8798 8678 8844 8730
rect 8844 8678 8854 8730
rect 8878 8678 8908 8730
rect 8908 8678 8920 8730
rect 8920 8678 8934 8730
rect 8958 8678 8972 8730
rect 8972 8678 8984 8730
rect 8984 8678 9014 8730
rect 9038 8678 9048 8730
rect 9048 8678 9094 8730
rect 8798 8676 8854 8678
rect 8878 8676 8934 8678
rect 8958 8676 9014 8678
rect 9038 8676 9094 8678
rect 16640 8730 16696 8732
rect 16720 8730 16776 8732
rect 16800 8730 16856 8732
rect 16880 8730 16936 8732
rect 16640 8678 16686 8730
rect 16686 8678 16696 8730
rect 16720 8678 16750 8730
rect 16750 8678 16762 8730
rect 16762 8678 16776 8730
rect 16800 8678 16814 8730
rect 16814 8678 16826 8730
rect 16826 8678 16856 8730
rect 16880 8678 16890 8730
rect 16890 8678 16936 8730
rect 16640 8676 16696 8678
rect 16720 8676 16776 8678
rect 16800 8676 16856 8678
rect 16880 8676 16936 8678
rect 24482 8730 24538 8732
rect 24562 8730 24618 8732
rect 24642 8730 24698 8732
rect 24722 8730 24778 8732
rect 24482 8678 24528 8730
rect 24528 8678 24538 8730
rect 24562 8678 24592 8730
rect 24592 8678 24604 8730
rect 24604 8678 24618 8730
rect 24642 8678 24656 8730
rect 24656 8678 24668 8730
rect 24668 8678 24698 8730
rect 24722 8678 24732 8730
rect 24732 8678 24778 8730
rect 24482 8676 24538 8678
rect 24562 8676 24618 8678
rect 24642 8676 24698 8678
rect 24722 8676 24778 8678
rect 32324 8730 32380 8732
rect 32404 8730 32460 8732
rect 32484 8730 32540 8732
rect 32564 8730 32620 8732
rect 32324 8678 32370 8730
rect 32370 8678 32380 8730
rect 32404 8678 32434 8730
rect 32434 8678 32446 8730
rect 32446 8678 32460 8730
rect 32484 8678 32498 8730
rect 32498 8678 32510 8730
rect 32510 8678 32540 8730
rect 32564 8678 32574 8730
rect 32574 8678 32620 8730
rect 32324 8676 32380 8678
rect 32404 8676 32460 8678
rect 32484 8676 32540 8678
rect 32564 8676 32620 8678
rect 4877 8186 4933 8188
rect 4957 8186 5013 8188
rect 5037 8186 5093 8188
rect 5117 8186 5173 8188
rect 4877 8134 4923 8186
rect 4923 8134 4933 8186
rect 4957 8134 4987 8186
rect 4987 8134 4999 8186
rect 4999 8134 5013 8186
rect 5037 8134 5051 8186
rect 5051 8134 5063 8186
rect 5063 8134 5093 8186
rect 5117 8134 5127 8186
rect 5127 8134 5173 8186
rect 4877 8132 4933 8134
rect 4957 8132 5013 8134
rect 5037 8132 5093 8134
rect 5117 8132 5173 8134
rect 12719 8186 12775 8188
rect 12799 8186 12855 8188
rect 12879 8186 12935 8188
rect 12959 8186 13015 8188
rect 12719 8134 12765 8186
rect 12765 8134 12775 8186
rect 12799 8134 12829 8186
rect 12829 8134 12841 8186
rect 12841 8134 12855 8186
rect 12879 8134 12893 8186
rect 12893 8134 12905 8186
rect 12905 8134 12935 8186
rect 12959 8134 12969 8186
rect 12969 8134 13015 8186
rect 12719 8132 12775 8134
rect 12799 8132 12855 8134
rect 12879 8132 12935 8134
rect 12959 8132 13015 8134
rect 20561 8186 20617 8188
rect 20641 8186 20697 8188
rect 20721 8186 20777 8188
rect 20801 8186 20857 8188
rect 20561 8134 20607 8186
rect 20607 8134 20617 8186
rect 20641 8134 20671 8186
rect 20671 8134 20683 8186
rect 20683 8134 20697 8186
rect 20721 8134 20735 8186
rect 20735 8134 20747 8186
rect 20747 8134 20777 8186
rect 20801 8134 20811 8186
rect 20811 8134 20857 8186
rect 20561 8132 20617 8134
rect 20641 8132 20697 8134
rect 20721 8132 20777 8134
rect 20801 8132 20857 8134
rect 28403 8186 28459 8188
rect 28483 8186 28539 8188
rect 28563 8186 28619 8188
rect 28643 8186 28699 8188
rect 28403 8134 28449 8186
rect 28449 8134 28459 8186
rect 28483 8134 28513 8186
rect 28513 8134 28525 8186
rect 28525 8134 28539 8186
rect 28563 8134 28577 8186
rect 28577 8134 28589 8186
rect 28589 8134 28619 8186
rect 28643 8134 28653 8186
rect 28653 8134 28699 8186
rect 28403 8132 28459 8134
rect 28483 8132 28539 8134
rect 28563 8132 28619 8134
rect 28643 8132 28699 8134
rect 8798 7642 8854 7644
rect 8878 7642 8934 7644
rect 8958 7642 9014 7644
rect 9038 7642 9094 7644
rect 8798 7590 8844 7642
rect 8844 7590 8854 7642
rect 8878 7590 8908 7642
rect 8908 7590 8920 7642
rect 8920 7590 8934 7642
rect 8958 7590 8972 7642
rect 8972 7590 8984 7642
rect 8984 7590 9014 7642
rect 9038 7590 9048 7642
rect 9048 7590 9094 7642
rect 8798 7588 8854 7590
rect 8878 7588 8934 7590
rect 8958 7588 9014 7590
rect 9038 7588 9094 7590
rect 16640 7642 16696 7644
rect 16720 7642 16776 7644
rect 16800 7642 16856 7644
rect 16880 7642 16936 7644
rect 16640 7590 16686 7642
rect 16686 7590 16696 7642
rect 16720 7590 16750 7642
rect 16750 7590 16762 7642
rect 16762 7590 16776 7642
rect 16800 7590 16814 7642
rect 16814 7590 16826 7642
rect 16826 7590 16856 7642
rect 16880 7590 16890 7642
rect 16890 7590 16936 7642
rect 16640 7588 16696 7590
rect 16720 7588 16776 7590
rect 16800 7588 16856 7590
rect 16880 7588 16936 7590
rect 24482 7642 24538 7644
rect 24562 7642 24618 7644
rect 24642 7642 24698 7644
rect 24722 7642 24778 7644
rect 24482 7590 24528 7642
rect 24528 7590 24538 7642
rect 24562 7590 24592 7642
rect 24592 7590 24604 7642
rect 24604 7590 24618 7642
rect 24642 7590 24656 7642
rect 24656 7590 24668 7642
rect 24668 7590 24698 7642
rect 24722 7590 24732 7642
rect 24732 7590 24778 7642
rect 24482 7588 24538 7590
rect 24562 7588 24618 7590
rect 24642 7588 24698 7590
rect 24722 7588 24778 7590
rect 32324 7642 32380 7644
rect 32404 7642 32460 7644
rect 32484 7642 32540 7644
rect 32564 7642 32620 7644
rect 32324 7590 32370 7642
rect 32370 7590 32380 7642
rect 32404 7590 32434 7642
rect 32434 7590 32446 7642
rect 32446 7590 32460 7642
rect 32484 7590 32498 7642
rect 32498 7590 32510 7642
rect 32510 7590 32540 7642
rect 32564 7590 32574 7642
rect 32574 7590 32620 7642
rect 32324 7588 32380 7590
rect 32404 7588 32460 7590
rect 32484 7588 32540 7590
rect 32564 7588 32620 7590
rect 4877 7098 4933 7100
rect 4957 7098 5013 7100
rect 5037 7098 5093 7100
rect 5117 7098 5173 7100
rect 4877 7046 4923 7098
rect 4923 7046 4933 7098
rect 4957 7046 4987 7098
rect 4987 7046 4999 7098
rect 4999 7046 5013 7098
rect 5037 7046 5051 7098
rect 5051 7046 5063 7098
rect 5063 7046 5093 7098
rect 5117 7046 5127 7098
rect 5127 7046 5173 7098
rect 4877 7044 4933 7046
rect 4957 7044 5013 7046
rect 5037 7044 5093 7046
rect 5117 7044 5173 7046
rect 12719 7098 12775 7100
rect 12799 7098 12855 7100
rect 12879 7098 12935 7100
rect 12959 7098 13015 7100
rect 12719 7046 12765 7098
rect 12765 7046 12775 7098
rect 12799 7046 12829 7098
rect 12829 7046 12841 7098
rect 12841 7046 12855 7098
rect 12879 7046 12893 7098
rect 12893 7046 12905 7098
rect 12905 7046 12935 7098
rect 12959 7046 12969 7098
rect 12969 7046 13015 7098
rect 12719 7044 12775 7046
rect 12799 7044 12855 7046
rect 12879 7044 12935 7046
rect 12959 7044 13015 7046
rect 20561 7098 20617 7100
rect 20641 7098 20697 7100
rect 20721 7098 20777 7100
rect 20801 7098 20857 7100
rect 20561 7046 20607 7098
rect 20607 7046 20617 7098
rect 20641 7046 20671 7098
rect 20671 7046 20683 7098
rect 20683 7046 20697 7098
rect 20721 7046 20735 7098
rect 20735 7046 20747 7098
rect 20747 7046 20777 7098
rect 20801 7046 20811 7098
rect 20811 7046 20857 7098
rect 20561 7044 20617 7046
rect 20641 7044 20697 7046
rect 20721 7044 20777 7046
rect 20801 7044 20857 7046
rect 28403 7098 28459 7100
rect 28483 7098 28539 7100
rect 28563 7098 28619 7100
rect 28643 7098 28699 7100
rect 28403 7046 28449 7098
rect 28449 7046 28459 7098
rect 28483 7046 28513 7098
rect 28513 7046 28525 7098
rect 28525 7046 28539 7098
rect 28563 7046 28577 7098
rect 28577 7046 28589 7098
rect 28589 7046 28619 7098
rect 28643 7046 28653 7098
rect 28653 7046 28699 7098
rect 28403 7044 28459 7046
rect 28483 7044 28539 7046
rect 28563 7044 28619 7046
rect 28643 7044 28699 7046
rect 8798 6554 8854 6556
rect 8878 6554 8934 6556
rect 8958 6554 9014 6556
rect 9038 6554 9094 6556
rect 8798 6502 8844 6554
rect 8844 6502 8854 6554
rect 8878 6502 8908 6554
rect 8908 6502 8920 6554
rect 8920 6502 8934 6554
rect 8958 6502 8972 6554
rect 8972 6502 8984 6554
rect 8984 6502 9014 6554
rect 9038 6502 9048 6554
rect 9048 6502 9094 6554
rect 8798 6500 8854 6502
rect 8878 6500 8934 6502
rect 8958 6500 9014 6502
rect 9038 6500 9094 6502
rect 16640 6554 16696 6556
rect 16720 6554 16776 6556
rect 16800 6554 16856 6556
rect 16880 6554 16936 6556
rect 16640 6502 16686 6554
rect 16686 6502 16696 6554
rect 16720 6502 16750 6554
rect 16750 6502 16762 6554
rect 16762 6502 16776 6554
rect 16800 6502 16814 6554
rect 16814 6502 16826 6554
rect 16826 6502 16856 6554
rect 16880 6502 16890 6554
rect 16890 6502 16936 6554
rect 16640 6500 16696 6502
rect 16720 6500 16776 6502
rect 16800 6500 16856 6502
rect 16880 6500 16936 6502
rect 24482 6554 24538 6556
rect 24562 6554 24618 6556
rect 24642 6554 24698 6556
rect 24722 6554 24778 6556
rect 24482 6502 24528 6554
rect 24528 6502 24538 6554
rect 24562 6502 24592 6554
rect 24592 6502 24604 6554
rect 24604 6502 24618 6554
rect 24642 6502 24656 6554
rect 24656 6502 24668 6554
rect 24668 6502 24698 6554
rect 24722 6502 24732 6554
rect 24732 6502 24778 6554
rect 24482 6500 24538 6502
rect 24562 6500 24618 6502
rect 24642 6500 24698 6502
rect 24722 6500 24778 6502
rect 32324 6554 32380 6556
rect 32404 6554 32460 6556
rect 32484 6554 32540 6556
rect 32564 6554 32620 6556
rect 32324 6502 32370 6554
rect 32370 6502 32380 6554
rect 32404 6502 32434 6554
rect 32434 6502 32446 6554
rect 32446 6502 32460 6554
rect 32484 6502 32498 6554
rect 32498 6502 32510 6554
rect 32510 6502 32540 6554
rect 32564 6502 32574 6554
rect 32574 6502 32620 6554
rect 32324 6500 32380 6502
rect 32404 6500 32460 6502
rect 32484 6500 32540 6502
rect 32564 6500 32620 6502
rect 4877 6010 4933 6012
rect 4957 6010 5013 6012
rect 5037 6010 5093 6012
rect 5117 6010 5173 6012
rect 4877 5958 4923 6010
rect 4923 5958 4933 6010
rect 4957 5958 4987 6010
rect 4987 5958 4999 6010
rect 4999 5958 5013 6010
rect 5037 5958 5051 6010
rect 5051 5958 5063 6010
rect 5063 5958 5093 6010
rect 5117 5958 5127 6010
rect 5127 5958 5173 6010
rect 4877 5956 4933 5958
rect 4957 5956 5013 5958
rect 5037 5956 5093 5958
rect 5117 5956 5173 5958
rect 12719 6010 12775 6012
rect 12799 6010 12855 6012
rect 12879 6010 12935 6012
rect 12959 6010 13015 6012
rect 12719 5958 12765 6010
rect 12765 5958 12775 6010
rect 12799 5958 12829 6010
rect 12829 5958 12841 6010
rect 12841 5958 12855 6010
rect 12879 5958 12893 6010
rect 12893 5958 12905 6010
rect 12905 5958 12935 6010
rect 12959 5958 12969 6010
rect 12969 5958 13015 6010
rect 12719 5956 12775 5958
rect 12799 5956 12855 5958
rect 12879 5956 12935 5958
rect 12959 5956 13015 5958
rect 20561 6010 20617 6012
rect 20641 6010 20697 6012
rect 20721 6010 20777 6012
rect 20801 6010 20857 6012
rect 20561 5958 20607 6010
rect 20607 5958 20617 6010
rect 20641 5958 20671 6010
rect 20671 5958 20683 6010
rect 20683 5958 20697 6010
rect 20721 5958 20735 6010
rect 20735 5958 20747 6010
rect 20747 5958 20777 6010
rect 20801 5958 20811 6010
rect 20811 5958 20857 6010
rect 20561 5956 20617 5958
rect 20641 5956 20697 5958
rect 20721 5956 20777 5958
rect 20801 5956 20857 5958
rect 28403 6010 28459 6012
rect 28483 6010 28539 6012
rect 28563 6010 28619 6012
rect 28643 6010 28699 6012
rect 28403 5958 28449 6010
rect 28449 5958 28459 6010
rect 28483 5958 28513 6010
rect 28513 5958 28525 6010
rect 28525 5958 28539 6010
rect 28563 5958 28577 6010
rect 28577 5958 28589 6010
rect 28589 5958 28619 6010
rect 28643 5958 28653 6010
rect 28653 5958 28699 6010
rect 28403 5956 28459 5958
rect 28483 5956 28539 5958
rect 28563 5956 28619 5958
rect 28643 5956 28699 5958
rect 8798 5466 8854 5468
rect 8878 5466 8934 5468
rect 8958 5466 9014 5468
rect 9038 5466 9094 5468
rect 8798 5414 8844 5466
rect 8844 5414 8854 5466
rect 8878 5414 8908 5466
rect 8908 5414 8920 5466
rect 8920 5414 8934 5466
rect 8958 5414 8972 5466
rect 8972 5414 8984 5466
rect 8984 5414 9014 5466
rect 9038 5414 9048 5466
rect 9048 5414 9094 5466
rect 8798 5412 8854 5414
rect 8878 5412 8934 5414
rect 8958 5412 9014 5414
rect 9038 5412 9094 5414
rect 16640 5466 16696 5468
rect 16720 5466 16776 5468
rect 16800 5466 16856 5468
rect 16880 5466 16936 5468
rect 16640 5414 16686 5466
rect 16686 5414 16696 5466
rect 16720 5414 16750 5466
rect 16750 5414 16762 5466
rect 16762 5414 16776 5466
rect 16800 5414 16814 5466
rect 16814 5414 16826 5466
rect 16826 5414 16856 5466
rect 16880 5414 16890 5466
rect 16890 5414 16936 5466
rect 16640 5412 16696 5414
rect 16720 5412 16776 5414
rect 16800 5412 16856 5414
rect 16880 5412 16936 5414
rect 24482 5466 24538 5468
rect 24562 5466 24618 5468
rect 24642 5466 24698 5468
rect 24722 5466 24778 5468
rect 24482 5414 24528 5466
rect 24528 5414 24538 5466
rect 24562 5414 24592 5466
rect 24592 5414 24604 5466
rect 24604 5414 24618 5466
rect 24642 5414 24656 5466
rect 24656 5414 24668 5466
rect 24668 5414 24698 5466
rect 24722 5414 24732 5466
rect 24732 5414 24778 5466
rect 24482 5412 24538 5414
rect 24562 5412 24618 5414
rect 24642 5412 24698 5414
rect 24722 5412 24778 5414
rect 32324 5466 32380 5468
rect 32404 5466 32460 5468
rect 32484 5466 32540 5468
rect 32564 5466 32620 5468
rect 32324 5414 32370 5466
rect 32370 5414 32380 5466
rect 32404 5414 32434 5466
rect 32434 5414 32446 5466
rect 32446 5414 32460 5466
rect 32484 5414 32498 5466
rect 32498 5414 32510 5466
rect 32510 5414 32540 5466
rect 32564 5414 32574 5466
rect 32574 5414 32620 5466
rect 32324 5412 32380 5414
rect 32404 5412 32460 5414
rect 32484 5412 32540 5414
rect 32564 5412 32620 5414
rect 4877 4922 4933 4924
rect 4957 4922 5013 4924
rect 5037 4922 5093 4924
rect 5117 4922 5173 4924
rect 4877 4870 4923 4922
rect 4923 4870 4933 4922
rect 4957 4870 4987 4922
rect 4987 4870 4999 4922
rect 4999 4870 5013 4922
rect 5037 4870 5051 4922
rect 5051 4870 5063 4922
rect 5063 4870 5093 4922
rect 5117 4870 5127 4922
rect 5127 4870 5173 4922
rect 4877 4868 4933 4870
rect 4957 4868 5013 4870
rect 5037 4868 5093 4870
rect 5117 4868 5173 4870
rect 12719 4922 12775 4924
rect 12799 4922 12855 4924
rect 12879 4922 12935 4924
rect 12959 4922 13015 4924
rect 12719 4870 12765 4922
rect 12765 4870 12775 4922
rect 12799 4870 12829 4922
rect 12829 4870 12841 4922
rect 12841 4870 12855 4922
rect 12879 4870 12893 4922
rect 12893 4870 12905 4922
rect 12905 4870 12935 4922
rect 12959 4870 12969 4922
rect 12969 4870 13015 4922
rect 12719 4868 12775 4870
rect 12799 4868 12855 4870
rect 12879 4868 12935 4870
rect 12959 4868 13015 4870
rect 20561 4922 20617 4924
rect 20641 4922 20697 4924
rect 20721 4922 20777 4924
rect 20801 4922 20857 4924
rect 20561 4870 20607 4922
rect 20607 4870 20617 4922
rect 20641 4870 20671 4922
rect 20671 4870 20683 4922
rect 20683 4870 20697 4922
rect 20721 4870 20735 4922
rect 20735 4870 20747 4922
rect 20747 4870 20777 4922
rect 20801 4870 20811 4922
rect 20811 4870 20857 4922
rect 20561 4868 20617 4870
rect 20641 4868 20697 4870
rect 20721 4868 20777 4870
rect 20801 4868 20857 4870
rect 28403 4922 28459 4924
rect 28483 4922 28539 4924
rect 28563 4922 28619 4924
rect 28643 4922 28699 4924
rect 28403 4870 28449 4922
rect 28449 4870 28459 4922
rect 28483 4870 28513 4922
rect 28513 4870 28525 4922
rect 28525 4870 28539 4922
rect 28563 4870 28577 4922
rect 28577 4870 28589 4922
rect 28589 4870 28619 4922
rect 28643 4870 28653 4922
rect 28653 4870 28699 4922
rect 28403 4868 28459 4870
rect 28483 4868 28539 4870
rect 28563 4868 28619 4870
rect 28643 4868 28699 4870
rect 8798 4378 8854 4380
rect 8878 4378 8934 4380
rect 8958 4378 9014 4380
rect 9038 4378 9094 4380
rect 8798 4326 8844 4378
rect 8844 4326 8854 4378
rect 8878 4326 8908 4378
rect 8908 4326 8920 4378
rect 8920 4326 8934 4378
rect 8958 4326 8972 4378
rect 8972 4326 8984 4378
rect 8984 4326 9014 4378
rect 9038 4326 9048 4378
rect 9048 4326 9094 4378
rect 8798 4324 8854 4326
rect 8878 4324 8934 4326
rect 8958 4324 9014 4326
rect 9038 4324 9094 4326
rect 16640 4378 16696 4380
rect 16720 4378 16776 4380
rect 16800 4378 16856 4380
rect 16880 4378 16936 4380
rect 16640 4326 16686 4378
rect 16686 4326 16696 4378
rect 16720 4326 16750 4378
rect 16750 4326 16762 4378
rect 16762 4326 16776 4378
rect 16800 4326 16814 4378
rect 16814 4326 16826 4378
rect 16826 4326 16856 4378
rect 16880 4326 16890 4378
rect 16890 4326 16936 4378
rect 16640 4324 16696 4326
rect 16720 4324 16776 4326
rect 16800 4324 16856 4326
rect 16880 4324 16936 4326
rect 24482 4378 24538 4380
rect 24562 4378 24618 4380
rect 24642 4378 24698 4380
rect 24722 4378 24778 4380
rect 24482 4326 24528 4378
rect 24528 4326 24538 4378
rect 24562 4326 24592 4378
rect 24592 4326 24604 4378
rect 24604 4326 24618 4378
rect 24642 4326 24656 4378
rect 24656 4326 24668 4378
rect 24668 4326 24698 4378
rect 24722 4326 24732 4378
rect 24732 4326 24778 4378
rect 24482 4324 24538 4326
rect 24562 4324 24618 4326
rect 24642 4324 24698 4326
rect 24722 4324 24778 4326
rect 32324 4378 32380 4380
rect 32404 4378 32460 4380
rect 32484 4378 32540 4380
rect 32564 4378 32620 4380
rect 32324 4326 32370 4378
rect 32370 4326 32380 4378
rect 32404 4326 32434 4378
rect 32434 4326 32446 4378
rect 32446 4326 32460 4378
rect 32484 4326 32498 4378
rect 32498 4326 32510 4378
rect 32510 4326 32540 4378
rect 32564 4326 32574 4378
rect 32574 4326 32620 4378
rect 32324 4324 32380 4326
rect 32404 4324 32460 4326
rect 32484 4324 32540 4326
rect 32564 4324 32620 4326
rect 4877 3834 4933 3836
rect 4957 3834 5013 3836
rect 5037 3834 5093 3836
rect 5117 3834 5173 3836
rect 4877 3782 4923 3834
rect 4923 3782 4933 3834
rect 4957 3782 4987 3834
rect 4987 3782 4999 3834
rect 4999 3782 5013 3834
rect 5037 3782 5051 3834
rect 5051 3782 5063 3834
rect 5063 3782 5093 3834
rect 5117 3782 5127 3834
rect 5127 3782 5173 3834
rect 4877 3780 4933 3782
rect 4957 3780 5013 3782
rect 5037 3780 5093 3782
rect 5117 3780 5173 3782
rect 12719 3834 12775 3836
rect 12799 3834 12855 3836
rect 12879 3834 12935 3836
rect 12959 3834 13015 3836
rect 12719 3782 12765 3834
rect 12765 3782 12775 3834
rect 12799 3782 12829 3834
rect 12829 3782 12841 3834
rect 12841 3782 12855 3834
rect 12879 3782 12893 3834
rect 12893 3782 12905 3834
rect 12905 3782 12935 3834
rect 12959 3782 12969 3834
rect 12969 3782 13015 3834
rect 12719 3780 12775 3782
rect 12799 3780 12855 3782
rect 12879 3780 12935 3782
rect 12959 3780 13015 3782
rect 20561 3834 20617 3836
rect 20641 3834 20697 3836
rect 20721 3834 20777 3836
rect 20801 3834 20857 3836
rect 20561 3782 20607 3834
rect 20607 3782 20617 3834
rect 20641 3782 20671 3834
rect 20671 3782 20683 3834
rect 20683 3782 20697 3834
rect 20721 3782 20735 3834
rect 20735 3782 20747 3834
rect 20747 3782 20777 3834
rect 20801 3782 20811 3834
rect 20811 3782 20857 3834
rect 20561 3780 20617 3782
rect 20641 3780 20697 3782
rect 20721 3780 20777 3782
rect 20801 3780 20857 3782
rect 28403 3834 28459 3836
rect 28483 3834 28539 3836
rect 28563 3834 28619 3836
rect 28643 3834 28699 3836
rect 28403 3782 28449 3834
rect 28449 3782 28459 3834
rect 28483 3782 28513 3834
rect 28513 3782 28525 3834
rect 28525 3782 28539 3834
rect 28563 3782 28577 3834
rect 28577 3782 28589 3834
rect 28589 3782 28619 3834
rect 28643 3782 28653 3834
rect 28653 3782 28699 3834
rect 28403 3780 28459 3782
rect 28483 3780 28539 3782
rect 28563 3780 28619 3782
rect 28643 3780 28699 3782
rect 8798 3290 8854 3292
rect 8878 3290 8934 3292
rect 8958 3290 9014 3292
rect 9038 3290 9094 3292
rect 8798 3238 8844 3290
rect 8844 3238 8854 3290
rect 8878 3238 8908 3290
rect 8908 3238 8920 3290
rect 8920 3238 8934 3290
rect 8958 3238 8972 3290
rect 8972 3238 8984 3290
rect 8984 3238 9014 3290
rect 9038 3238 9048 3290
rect 9048 3238 9094 3290
rect 8798 3236 8854 3238
rect 8878 3236 8934 3238
rect 8958 3236 9014 3238
rect 9038 3236 9094 3238
rect 16640 3290 16696 3292
rect 16720 3290 16776 3292
rect 16800 3290 16856 3292
rect 16880 3290 16936 3292
rect 16640 3238 16686 3290
rect 16686 3238 16696 3290
rect 16720 3238 16750 3290
rect 16750 3238 16762 3290
rect 16762 3238 16776 3290
rect 16800 3238 16814 3290
rect 16814 3238 16826 3290
rect 16826 3238 16856 3290
rect 16880 3238 16890 3290
rect 16890 3238 16936 3290
rect 16640 3236 16696 3238
rect 16720 3236 16776 3238
rect 16800 3236 16856 3238
rect 16880 3236 16936 3238
rect 24482 3290 24538 3292
rect 24562 3290 24618 3292
rect 24642 3290 24698 3292
rect 24722 3290 24778 3292
rect 24482 3238 24528 3290
rect 24528 3238 24538 3290
rect 24562 3238 24592 3290
rect 24592 3238 24604 3290
rect 24604 3238 24618 3290
rect 24642 3238 24656 3290
rect 24656 3238 24668 3290
rect 24668 3238 24698 3290
rect 24722 3238 24732 3290
rect 24732 3238 24778 3290
rect 24482 3236 24538 3238
rect 24562 3236 24618 3238
rect 24642 3236 24698 3238
rect 24722 3236 24778 3238
rect 32324 3290 32380 3292
rect 32404 3290 32460 3292
rect 32484 3290 32540 3292
rect 32564 3290 32620 3292
rect 32324 3238 32370 3290
rect 32370 3238 32380 3290
rect 32404 3238 32434 3290
rect 32434 3238 32446 3290
rect 32446 3238 32460 3290
rect 32484 3238 32498 3290
rect 32498 3238 32510 3290
rect 32510 3238 32540 3290
rect 32564 3238 32574 3290
rect 32574 3238 32620 3290
rect 32324 3236 32380 3238
rect 32404 3236 32460 3238
rect 32484 3236 32540 3238
rect 32564 3236 32620 3238
rect 4877 2746 4933 2748
rect 4957 2746 5013 2748
rect 5037 2746 5093 2748
rect 5117 2746 5173 2748
rect 4877 2694 4923 2746
rect 4923 2694 4933 2746
rect 4957 2694 4987 2746
rect 4987 2694 4999 2746
rect 4999 2694 5013 2746
rect 5037 2694 5051 2746
rect 5051 2694 5063 2746
rect 5063 2694 5093 2746
rect 5117 2694 5127 2746
rect 5127 2694 5173 2746
rect 4877 2692 4933 2694
rect 4957 2692 5013 2694
rect 5037 2692 5093 2694
rect 5117 2692 5173 2694
rect 12719 2746 12775 2748
rect 12799 2746 12855 2748
rect 12879 2746 12935 2748
rect 12959 2746 13015 2748
rect 12719 2694 12765 2746
rect 12765 2694 12775 2746
rect 12799 2694 12829 2746
rect 12829 2694 12841 2746
rect 12841 2694 12855 2746
rect 12879 2694 12893 2746
rect 12893 2694 12905 2746
rect 12905 2694 12935 2746
rect 12959 2694 12969 2746
rect 12969 2694 13015 2746
rect 12719 2692 12775 2694
rect 12799 2692 12855 2694
rect 12879 2692 12935 2694
rect 12959 2692 13015 2694
rect 20561 2746 20617 2748
rect 20641 2746 20697 2748
rect 20721 2746 20777 2748
rect 20801 2746 20857 2748
rect 20561 2694 20607 2746
rect 20607 2694 20617 2746
rect 20641 2694 20671 2746
rect 20671 2694 20683 2746
rect 20683 2694 20697 2746
rect 20721 2694 20735 2746
rect 20735 2694 20747 2746
rect 20747 2694 20777 2746
rect 20801 2694 20811 2746
rect 20811 2694 20857 2746
rect 20561 2692 20617 2694
rect 20641 2692 20697 2694
rect 20721 2692 20777 2694
rect 20801 2692 20857 2694
rect 28403 2746 28459 2748
rect 28483 2746 28539 2748
rect 28563 2746 28619 2748
rect 28643 2746 28699 2748
rect 28403 2694 28449 2746
rect 28449 2694 28459 2746
rect 28483 2694 28513 2746
rect 28513 2694 28525 2746
rect 28525 2694 28539 2746
rect 28563 2694 28577 2746
rect 28577 2694 28589 2746
rect 28589 2694 28619 2746
rect 28643 2694 28653 2746
rect 28653 2694 28699 2746
rect 28403 2692 28459 2694
rect 28483 2692 28539 2694
rect 28563 2692 28619 2694
rect 28643 2692 28699 2694
rect 8798 2202 8854 2204
rect 8878 2202 8934 2204
rect 8958 2202 9014 2204
rect 9038 2202 9094 2204
rect 8798 2150 8844 2202
rect 8844 2150 8854 2202
rect 8878 2150 8908 2202
rect 8908 2150 8920 2202
rect 8920 2150 8934 2202
rect 8958 2150 8972 2202
rect 8972 2150 8984 2202
rect 8984 2150 9014 2202
rect 9038 2150 9048 2202
rect 9048 2150 9094 2202
rect 8798 2148 8854 2150
rect 8878 2148 8934 2150
rect 8958 2148 9014 2150
rect 9038 2148 9094 2150
rect 16640 2202 16696 2204
rect 16720 2202 16776 2204
rect 16800 2202 16856 2204
rect 16880 2202 16936 2204
rect 16640 2150 16686 2202
rect 16686 2150 16696 2202
rect 16720 2150 16750 2202
rect 16750 2150 16762 2202
rect 16762 2150 16776 2202
rect 16800 2150 16814 2202
rect 16814 2150 16826 2202
rect 16826 2150 16856 2202
rect 16880 2150 16890 2202
rect 16890 2150 16936 2202
rect 16640 2148 16696 2150
rect 16720 2148 16776 2150
rect 16800 2148 16856 2150
rect 16880 2148 16936 2150
rect 24482 2202 24538 2204
rect 24562 2202 24618 2204
rect 24642 2202 24698 2204
rect 24722 2202 24778 2204
rect 24482 2150 24528 2202
rect 24528 2150 24538 2202
rect 24562 2150 24592 2202
rect 24592 2150 24604 2202
rect 24604 2150 24618 2202
rect 24642 2150 24656 2202
rect 24656 2150 24668 2202
rect 24668 2150 24698 2202
rect 24722 2150 24732 2202
rect 24732 2150 24778 2202
rect 24482 2148 24538 2150
rect 24562 2148 24618 2150
rect 24642 2148 24698 2150
rect 24722 2148 24778 2150
rect 32324 2202 32380 2204
rect 32404 2202 32460 2204
rect 32484 2202 32540 2204
rect 32564 2202 32620 2204
rect 32324 2150 32370 2202
rect 32370 2150 32380 2202
rect 32404 2150 32434 2202
rect 32434 2150 32446 2202
rect 32446 2150 32460 2202
rect 32484 2150 32498 2202
rect 32498 2150 32510 2202
rect 32510 2150 32540 2202
rect 32564 2150 32574 2202
rect 32574 2150 32620 2202
rect 32324 2148 32380 2150
rect 32404 2148 32460 2150
rect 32484 2148 32540 2150
rect 32564 2148 32620 2150
rect 4877 1658 4933 1660
rect 4957 1658 5013 1660
rect 5037 1658 5093 1660
rect 5117 1658 5173 1660
rect 4877 1606 4923 1658
rect 4923 1606 4933 1658
rect 4957 1606 4987 1658
rect 4987 1606 4999 1658
rect 4999 1606 5013 1658
rect 5037 1606 5051 1658
rect 5051 1606 5063 1658
rect 5063 1606 5093 1658
rect 5117 1606 5127 1658
rect 5127 1606 5173 1658
rect 4877 1604 4933 1606
rect 4957 1604 5013 1606
rect 5037 1604 5093 1606
rect 5117 1604 5173 1606
rect 12719 1658 12775 1660
rect 12799 1658 12855 1660
rect 12879 1658 12935 1660
rect 12959 1658 13015 1660
rect 12719 1606 12765 1658
rect 12765 1606 12775 1658
rect 12799 1606 12829 1658
rect 12829 1606 12841 1658
rect 12841 1606 12855 1658
rect 12879 1606 12893 1658
rect 12893 1606 12905 1658
rect 12905 1606 12935 1658
rect 12959 1606 12969 1658
rect 12969 1606 13015 1658
rect 12719 1604 12775 1606
rect 12799 1604 12855 1606
rect 12879 1604 12935 1606
rect 12959 1604 13015 1606
rect 20561 1658 20617 1660
rect 20641 1658 20697 1660
rect 20721 1658 20777 1660
rect 20801 1658 20857 1660
rect 20561 1606 20607 1658
rect 20607 1606 20617 1658
rect 20641 1606 20671 1658
rect 20671 1606 20683 1658
rect 20683 1606 20697 1658
rect 20721 1606 20735 1658
rect 20735 1606 20747 1658
rect 20747 1606 20777 1658
rect 20801 1606 20811 1658
rect 20811 1606 20857 1658
rect 20561 1604 20617 1606
rect 20641 1604 20697 1606
rect 20721 1604 20777 1606
rect 20801 1604 20857 1606
rect 28403 1658 28459 1660
rect 28483 1658 28539 1660
rect 28563 1658 28619 1660
rect 28643 1658 28699 1660
rect 28403 1606 28449 1658
rect 28449 1606 28459 1658
rect 28483 1606 28513 1658
rect 28513 1606 28525 1658
rect 28525 1606 28539 1658
rect 28563 1606 28577 1658
rect 28577 1606 28589 1658
rect 28589 1606 28619 1658
rect 28643 1606 28653 1658
rect 28653 1606 28699 1658
rect 28403 1604 28459 1606
rect 28483 1604 28539 1606
rect 28563 1604 28619 1606
rect 28643 1604 28699 1606
rect 8798 1114 8854 1116
rect 8878 1114 8934 1116
rect 8958 1114 9014 1116
rect 9038 1114 9094 1116
rect 8798 1062 8844 1114
rect 8844 1062 8854 1114
rect 8878 1062 8908 1114
rect 8908 1062 8920 1114
rect 8920 1062 8934 1114
rect 8958 1062 8972 1114
rect 8972 1062 8984 1114
rect 8984 1062 9014 1114
rect 9038 1062 9048 1114
rect 9048 1062 9094 1114
rect 8798 1060 8854 1062
rect 8878 1060 8934 1062
rect 8958 1060 9014 1062
rect 9038 1060 9094 1062
rect 16640 1114 16696 1116
rect 16720 1114 16776 1116
rect 16800 1114 16856 1116
rect 16880 1114 16936 1116
rect 16640 1062 16686 1114
rect 16686 1062 16696 1114
rect 16720 1062 16750 1114
rect 16750 1062 16762 1114
rect 16762 1062 16776 1114
rect 16800 1062 16814 1114
rect 16814 1062 16826 1114
rect 16826 1062 16856 1114
rect 16880 1062 16890 1114
rect 16890 1062 16936 1114
rect 16640 1060 16696 1062
rect 16720 1060 16776 1062
rect 16800 1060 16856 1062
rect 16880 1060 16936 1062
rect 24482 1114 24538 1116
rect 24562 1114 24618 1116
rect 24642 1114 24698 1116
rect 24722 1114 24778 1116
rect 24482 1062 24528 1114
rect 24528 1062 24538 1114
rect 24562 1062 24592 1114
rect 24592 1062 24604 1114
rect 24604 1062 24618 1114
rect 24642 1062 24656 1114
rect 24656 1062 24668 1114
rect 24668 1062 24698 1114
rect 24722 1062 24732 1114
rect 24732 1062 24778 1114
rect 24482 1060 24538 1062
rect 24562 1060 24618 1062
rect 24642 1060 24698 1062
rect 24722 1060 24778 1062
rect 32324 1114 32380 1116
rect 32404 1114 32460 1116
rect 32484 1114 32540 1116
rect 32564 1114 32620 1116
rect 32324 1062 32370 1114
rect 32370 1062 32380 1114
rect 32404 1062 32434 1114
rect 32434 1062 32446 1114
rect 32446 1062 32460 1114
rect 32484 1062 32498 1114
rect 32498 1062 32510 1114
rect 32510 1062 32540 1114
rect 32564 1062 32574 1114
rect 32574 1062 32620 1114
rect 32324 1060 32380 1062
rect 32404 1060 32460 1062
rect 32484 1060 32540 1062
rect 32564 1060 32620 1062
<< metal3 >>
rect 8886 21388 8892 21452
rect 8956 21450 8962 21452
rect 9121 21450 9187 21453
rect 9673 21452 9739 21453
rect 8956 21448 9187 21450
rect 8956 21392 9126 21448
rect 9182 21392 9187 21448
rect 8956 21390 9187 21392
rect 8956 21388 8962 21390
rect 9121 21387 9187 21390
rect 9622 21388 9628 21452
rect 9692 21450 9739 21452
rect 11053 21452 11119 21453
rect 11881 21452 11947 21453
rect 11053 21450 11100 21452
rect 9692 21448 9784 21450
rect 9734 21392 9784 21448
rect 9692 21390 9784 21392
rect 11008 21448 11100 21450
rect 11008 21392 11058 21448
rect 11008 21390 11100 21392
rect 9692 21388 9739 21390
rect 9673 21387 9739 21388
rect 11053 21388 11100 21390
rect 11164 21388 11170 21452
rect 11830 21388 11836 21452
rect 11900 21450 11947 21452
rect 12801 21450 12867 21453
rect 13302 21450 13308 21452
rect 11900 21448 11992 21450
rect 11942 21392 11992 21448
rect 11900 21390 11992 21392
rect 12801 21448 13308 21450
rect 12801 21392 12806 21448
rect 12862 21392 13308 21448
rect 12801 21390 13308 21392
rect 11900 21388 11947 21390
rect 11053 21387 11119 21388
rect 11881 21387 11947 21388
rect 12801 21387 12867 21390
rect 13302 21388 13308 21390
rect 13372 21388 13378 21452
rect 13997 21450 14063 21453
rect 15561 21452 15627 21453
rect 14774 21450 14780 21452
rect 13997 21448 14780 21450
rect 13997 21392 14002 21448
rect 14058 21392 14780 21448
rect 13997 21390 14780 21392
rect 13997 21387 14063 21390
rect 14774 21388 14780 21390
rect 14844 21388 14850 21452
rect 15510 21450 15516 21452
rect 15470 21390 15516 21450
rect 15580 21448 15627 21452
rect 15622 21392 15627 21448
rect 15510 21388 15516 21390
rect 15580 21388 15627 21392
rect 15561 21387 15627 21388
rect 15745 21450 15811 21453
rect 16246 21450 16252 21452
rect 15745 21448 16252 21450
rect 15745 21392 15750 21448
rect 15806 21392 16252 21448
rect 15745 21390 16252 21392
rect 15745 21387 15811 21390
rect 16246 21388 16252 21390
rect 16316 21388 16322 21452
rect 17493 21450 17559 21453
rect 17718 21450 17724 21452
rect 17493 21448 17724 21450
rect 17493 21392 17498 21448
rect 17554 21392 17724 21448
rect 17493 21390 17724 21392
rect 17493 21387 17559 21390
rect 17718 21388 17724 21390
rect 17788 21388 17794 21452
rect 18454 21388 18460 21452
rect 18524 21450 18530 21452
rect 19241 21450 19307 21453
rect 18524 21448 19307 21450
rect 18524 21392 19246 21448
rect 19302 21392 19307 21448
rect 18524 21390 19307 21392
rect 18524 21388 18530 21390
rect 19241 21387 19307 21390
rect 19517 21450 19583 21453
rect 19926 21450 19932 21452
rect 19517 21448 19932 21450
rect 19517 21392 19522 21448
rect 19578 21392 19932 21448
rect 19517 21390 19932 21392
rect 19517 21387 19583 21390
rect 19926 21388 19932 21390
rect 19996 21388 20002 21452
rect 21398 21388 21404 21452
rect 21468 21450 21474 21452
rect 21725 21450 21791 21453
rect 21468 21448 21791 21450
rect 21468 21392 21730 21448
rect 21786 21392 21791 21448
rect 21468 21390 21791 21392
rect 21468 21388 21474 21390
rect 21725 21387 21791 21390
rect 22134 21388 22140 21452
rect 22204 21450 22210 21452
rect 22921 21450 22987 21453
rect 23657 21452 23723 21453
rect 24393 21452 24459 21453
rect 25865 21452 25931 21453
rect 23606 21450 23612 21452
rect 22204 21448 22987 21450
rect 22204 21392 22926 21448
rect 22982 21392 22987 21448
rect 22204 21390 22987 21392
rect 23566 21390 23612 21450
rect 23676 21448 23723 21452
rect 24342 21450 24348 21452
rect 23718 21392 23723 21448
rect 22204 21388 22210 21390
rect 22921 21387 22987 21390
rect 23606 21388 23612 21390
rect 23676 21388 23723 21392
rect 24302 21390 24348 21450
rect 24412 21448 24459 21452
rect 25814 21450 25820 21452
rect 24454 21392 24459 21448
rect 24342 21388 24348 21390
rect 24412 21388 24459 21392
rect 25774 21390 25820 21450
rect 25884 21448 25931 21452
rect 25926 21392 25931 21448
rect 25814 21388 25820 21390
rect 25884 21388 25931 21392
rect 27286 21388 27292 21452
rect 27356 21450 27362 21452
rect 27429 21450 27495 21453
rect 28809 21452 28875 21453
rect 30281 21452 30347 21453
rect 28758 21450 28764 21452
rect 27356 21448 27495 21450
rect 27356 21392 27434 21448
rect 27490 21392 27495 21448
rect 27356 21390 27495 21392
rect 28718 21390 28764 21450
rect 28828 21448 28875 21452
rect 30230 21450 30236 21452
rect 28870 21392 28875 21448
rect 27356 21388 27362 21390
rect 23657 21387 23723 21388
rect 24393 21387 24459 21388
rect 25865 21387 25931 21388
rect 27429 21387 27495 21390
rect 28758 21388 28764 21390
rect 28828 21388 28875 21392
rect 30190 21390 30236 21450
rect 30300 21448 30347 21452
rect 30342 21392 30347 21448
rect 30230 21388 30236 21390
rect 30300 21388 30347 21392
rect 28809 21387 28875 21388
rect 30281 21387 30347 21388
rect 13813 21314 13879 21317
rect 14038 21314 14044 21316
rect 13813 21312 14044 21314
rect 13813 21256 13818 21312
rect 13874 21256 14044 21312
rect 13813 21254 14044 21256
rect 13813 21251 13879 21254
rect 14038 21252 14044 21254
rect 14108 21252 14114 21316
rect 16982 21252 16988 21316
rect 17052 21314 17058 21316
rect 17861 21314 17927 21317
rect 17052 21312 17927 21314
rect 17052 21256 17866 21312
rect 17922 21256 17927 21312
rect 17052 21254 17927 21256
rect 17052 21252 17058 21254
rect 17861 21251 17927 21254
rect 20300 21274 20386 21282
rect 21208 21276 21316 21296
rect 21208 21274 21226 21276
rect 20300 21272 21226 21274
rect 20300 21208 20310 21272
rect 20374 21216 21226 21272
rect 21296 21216 21316 21276
rect 20374 21214 21316 21216
rect 20374 21208 20386 21214
rect 20300 21198 20386 21208
rect 21208 21198 21316 21214
rect 33598 21280 33714 21294
rect 33598 21208 33614 21280
rect 33696 21208 33714 21280
rect 33598 21192 33714 21208
rect 26550 20980 26556 21044
rect 26620 21042 26626 21044
rect 27337 21042 27403 21045
rect 26620 21040 27403 21042
rect 26620 20984 27342 21040
rect 27398 20984 27403 21040
rect 26620 20982 27403 20984
rect 26620 20980 26626 20982
rect 27337 20979 27403 20982
rect 28022 20980 28028 21044
rect 28092 21042 28098 21044
rect 28625 21042 28691 21045
rect 28092 21040 28691 21042
rect 28092 20984 28630 21040
rect 28686 20984 28691 21040
rect 28092 20982 28691 20984
rect 28092 20980 28098 20982
rect 28625 20979 28691 20982
rect 29494 20980 29500 21044
rect 29564 21042 29570 21044
rect 29913 21042 29979 21045
rect 29564 21040 29979 21042
rect 29564 20984 29918 21040
rect 29974 20984 29979 21040
rect 29564 20982 29979 20984
rect 29564 20980 29570 20982
rect 29913 20979 29979 20982
rect 5165 20908 5231 20909
rect 5165 20906 5212 20908
rect 5120 20904 5212 20906
rect 5120 20848 5170 20904
rect 5120 20846 5212 20848
rect 5165 20844 5212 20846
rect 5276 20844 5282 20908
rect 20662 20844 20668 20908
rect 20732 20906 20738 20908
rect 20897 20906 20963 20909
rect 20732 20904 20963 20906
rect 20732 20848 20902 20904
rect 20958 20848 20963 20904
rect 20732 20846 20963 20848
rect 20732 20844 20738 20846
rect 5165 20843 5231 20844
rect 20897 20843 20963 20846
rect 8788 20704 9104 20705
rect 8788 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8954 20704
rect 9018 20640 9034 20704
rect 9098 20640 9104 20704
rect 8788 20639 9104 20640
rect 16630 20704 16946 20705
rect 16630 20640 16636 20704
rect 16700 20640 16716 20704
rect 16780 20640 16796 20704
rect 16860 20640 16876 20704
rect 16940 20640 16946 20704
rect 16630 20639 16946 20640
rect 24472 20704 24788 20705
rect 24472 20640 24478 20704
rect 24542 20640 24558 20704
rect 24622 20640 24638 20704
rect 24702 20640 24718 20704
rect 24782 20640 24788 20704
rect 24472 20639 24788 20640
rect 32314 20704 32630 20705
rect 32314 20640 32320 20704
rect 32384 20640 32400 20704
rect 32464 20640 32480 20704
rect 32544 20640 32560 20704
rect 32624 20640 32630 20704
rect 32314 20639 32630 20640
rect 2129 20498 2195 20501
rect 2262 20498 2268 20500
rect 2129 20496 2268 20498
rect 2129 20440 2134 20496
rect 2190 20440 2268 20496
rect 2129 20438 2268 20440
rect 2129 20435 2195 20438
rect 2262 20436 2268 20438
rect 2332 20436 2338 20500
rect 2773 20498 2839 20501
rect 2998 20498 3004 20500
rect 2773 20496 3004 20498
rect 2773 20440 2778 20496
rect 2834 20440 3004 20496
rect 2773 20438 3004 20440
rect 2773 20435 2839 20438
rect 2998 20436 3004 20438
rect 3068 20436 3074 20500
rect 3417 20498 3483 20501
rect 4521 20500 4587 20501
rect 5993 20500 6059 20501
rect 3734 20498 3740 20500
rect 3417 20496 3740 20498
rect 3417 20440 3422 20496
rect 3478 20440 3740 20496
rect 3417 20438 3740 20440
rect 3417 20435 3483 20438
rect 3734 20436 3740 20438
rect 3804 20436 3810 20500
rect 4470 20436 4476 20500
rect 4540 20498 4587 20500
rect 4540 20496 4632 20498
rect 4582 20440 4632 20496
rect 4540 20438 4632 20440
rect 4540 20436 4587 20438
rect 5942 20436 5948 20500
rect 6012 20498 6059 20500
rect 6012 20496 6104 20498
rect 6054 20440 6104 20496
rect 6012 20438 6104 20440
rect 6012 20436 6059 20438
rect 22870 20436 22876 20500
rect 22940 20498 22946 20500
rect 24761 20498 24827 20501
rect 22940 20496 24827 20498
rect 22940 20440 24766 20496
rect 24822 20440 24827 20496
rect 22940 20438 24827 20440
rect 22940 20436 22946 20438
rect 4521 20435 4587 20436
rect 5993 20435 6059 20436
rect 24761 20435 24827 20438
rect 12617 20364 12683 20365
rect 12566 20300 12572 20364
rect 12636 20362 12683 20364
rect 12636 20360 12728 20362
rect 12678 20304 12728 20360
rect 12636 20302 12728 20304
rect 12636 20300 12683 20302
rect 12617 20299 12683 20300
rect 4867 20160 5183 20161
rect 4867 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5113 20160
rect 5177 20096 5183 20160
rect 4867 20095 5183 20096
rect 12709 20160 13025 20161
rect 12709 20096 12715 20160
rect 12779 20096 12795 20160
rect 12859 20096 12875 20160
rect 12939 20096 12955 20160
rect 13019 20096 13025 20160
rect 12709 20095 13025 20096
rect 20551 20160 20867 20161
rect 20551 20096 20557 20160
rect 20621 20096 20637 20160
rect 20701 20096 20717 20160
rect 20781 20096 20797 20160
rect 20861 20096 20867 20160
rect 20551 20095 20867 20096
rect 28393 20160 28709 20161
rect 28393 20096 28399 20160
rect 28463 20096 28479 20160
rect 28543 20096 28559 20160
rect 28623 20096 28639 20160
rect 28703 20096 28709 20160
rect 28393 20095 28709 20096
rect 1577 20092 1643 20093
rect 6729 20092 6795 20093
rect 7465 20092 7531 20093
rect 8201 20092 8267 20093
rect 1526 20028 1532 20092
rect 1596 20090 1643 20092
rect 1596 20088 1688 20090
rect 1638 20032 1688 20088
rect 1596 20030 1688 20032
rect 1596 20028 1643 20030
rect 6678 20028 6684 20092
rect 6748 20090 6795 20092
rect 6748 20088 6840 20090
rect 6790 20032 6840 20088
rect 6748 20030 6840 20032
rect 6748 20028 6795 20030
rect 7414 20028 7420 20092
rect 7484 20090 7531 20092
rect 7484 20088 7576 20090
rect 7526 20032 7576 20088
rect 7484 20030 7576 20032
rect 7484 20028 7531 20030
rect 8150 20028 8156 20092
rect 8220 20090 8267 20092
rect 10133 20090 10199 20093
rect 10358 20090 10364 20092
rect 8220 20088 8312 20090
rect 8262 20032 8312 20088
rect 8220 20030 8312 20032
rect 10133 20088 10364 20090
rect 10133 20032 10138 20088
rect 10194 20032 10364 20088
rect 10133 20030 10364 20032
rect 8220 20028 8267 20030
rect 1577 20027 1643 20028
rect 6729 20027 6795 20028
rect 7465 20027 7531 20028
rect 8201 20027 8267 20028
rect 10133 20027 10199 20030
rect 10358 20028 10364 20030
rect 10428 20028 10434 20092
rect 20805 19954 20871 19957
rect 21173 19954 21239 19957
rect 20805 19952 21239 19954
rect 20805 19896 20810 19952
rect 20866 19896 21178 19952
rect 21234 19896 21239 19952
rect 20805 19894 21239 19896
rect 20805 19891 20871 19894
rect 21173 19891 21239 19894
rect 8788 19616 9104 19617
rect 8788 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8954 19616
rect 9018 19552 9034 19616
rect 9098 19552 9104 19616
rect 8788 19551 9104 19552
rect 16630 19616 16946 19617
rect 16630 19552 16636 19616
rect 16700 19552 16716 19616
rect 16780 19552 16796 19616
rect 16860 19552 16876 19616
rect 16940 19552 16946 19616
rect 16630 19551 16946 19552
rect 24472 19616 24788 19617
rect 24472 19552 24478 19616
rect 24542 19552 24558 19616
rect 24622 19552 24638 19616
rect 24702 19552 24718 19616
rect 24782 19552 24788 19616
rect 24472 19551 24788 19552
rect 32314 19616 32630 19617
rect 32314 19552 32320 19616
rect 32384 19552 32400 19616
rect 32464 19552 32480 19616
rect 32544 19552 32560 19616
rect 32624 19552 32630 19616
rect 32314 19551 32630 19552
rect 21817 19546 21883 19549
rect 23565 19546 23631 19549
rect 21817 19544 23631 19546
rect 21817 19488 21822 19544
rect 21878 19488 23570 19544
rect 23626 19488 23631 19544
rect 21817 19486 23631 19488
rect 21817 19483 21883 19486
rect 23565 19483 23631 19486
rect 20621 19274 20687 19277
rect 22001 19274 22067 19277
rect 20621 19272 22067 19274
rect 20621 19216 20626 19272
rect 20682 19216 22006 19272
rect 22062 19216 22067 19272
rect 20621 19214 22067 19216
rect 20621 19211 20687 19214
rect 22001 19211 22067 19214
rect 4867 19072 5183 19073
rect 4867 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5113 19072
rect 5177 19008 5183 19072
rect 4867 19007 5183 19008
rect 12709 19072 13025 19073
rect 12709 19008 12715 19072
rect 12779 19008 12795 19072
rect 12859 19008 12875 19072
rect 12939 19008 12955 19072
rect 13019 19008 13025 19072
rect 12709 19007 13025 19008
rect 20551 19072 20867 19073
rect 20551 19008 20557 19072
rect 20621 19008 20637 19072
rect 20701 19008 20717 19072
rect 20781 19008 20797 19072
rect 20861 19008 20867 19072
rect 20551 19007 20867 19008
rect 28393 19072 28709 19073
rect 28393 19008 28399 19072
rect 28463 19008 28479 19072
rect 28543 19008 28559 19072
rect 28623 19008 28639 19072
rect 28703 19008 28709 19072
rect 28393 19007 28709 19008
rect 8788 18528 9104 18529
rect 8788 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8954 18528
rect 9018 18464 9034 18528
rect 9098 18464 9104 18528
rect 8788 18463 9104 18464
rect 16630 18528 16946 18529
rect 16630 18464 16636 18528
rect 16700 18464 16716 18528
rect 16780 18464 16796 18528
rect 16860 18464 16876 18528
rect 16940 18464 16946 18528
rect 16630 18463 16946 18464
rect 24472 18528 24788 18529
rect 24472 18464 24478 18528
rect 24542 18464 24558 18528
rect 24622 18464 24638 18528
rect 24702 18464 24718 18528
rect 24782 18464 24788 18528
rect 24472 18463 24788 18464
rect 32314 18528 32630 18529
rect 32314 18464 32320 18528
rect 32384 18464 32400 18528
rect 32464 18464 32480 18528
rect 32544 18464 32560 18528
rect 32624 18464 32630 18528
rect 32314 18463 32630 18464
rect 4867 17984 5183 17985
rect 4867 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5113 17984
rect 5177 17920 5183 17984
rect 4867 17919 5183 17920
rect 12709 17984 13025 17985
rect 12709 17920 12715 17984
rect 12779 17920 12795 17984
rect 12859 17920 12875 17984
rect 12939 17920 12955 17984
rect 13019 17920 13025 17984
rect 12709 17919 13025 17920
rect 20551 17984 20867 17985
rect 20551 17920 20557 17984
rect 20621 17920 20637 17984
rect 20701 17920 20717 17984
rect 20781 17920 20797 17984
rect 20861 17920 20867 17984
rect 20551 17919 20867 17920
rect 28393 17984 28709 17985
rect 28393 17920 28399 17984
rect 28463 17920 28479 17984
rect 28543 17920 28559 17984
rect 28623 17920 28639 17984
rect 28703 17920 28709 17984
rect 28393 17919 28709 17920
rect 8788 17440 9104 17441
rect 8788 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8954 17440
rect 9018 17376 9034 17440
rect 9098 17376 9104 17440
rect 8788 17375 9104 17376
rect 16630 17440 16946 17441
rect 16630 17376 16636 17440
rect 16700 17376 16716 17440
rect 16780 17376 16796 17440
rect 16860 17376 16876 17440
rect 16940 17376 16946 17440
rect 16630 17375 16946 17376
rect 24472 17440 24788 17441
rect 24472 17376 24478 17440
rect 24542 17376 24558 17440
rect 24622 17376 24638 17440
rect 24702 17376 24718 17440
rect 24782 17376 24788 17440
rect 24472 17375 24788 17376
rect 32314 17440 32630 17441
rect 32314 17376 32320 17440
rect 32384 17376 32400 17440
rect 32464 17376 32480 17440
rect 32544 17376 32560 17440
rect 32624 17376 32630 17440
rect 32314 17375 32630 17376
rect 4867 16896 5183 16897
rect 4867 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5113 16896
rect 5177 16832 5183 16896
rect 4867 16831 5183 16832
rect 12709 16896 13025 16897
rect 12709 16832 12715 16896
rect 12779 16832 12795 16896
rect 12859 16832 12875 16896
rect 12939 16832 12955 16896
rect 13019 16832 13025 16896
rect 12709 16831 13025 16832
rect 20551 16896 20867 16897
rect 20551 16832 20557 16896
rect 20621 16832 20637 16896
rect 20701 16832 20717 16896
rect 20781 16832 20797 16896
rect 20861 16832 20867 16896
rect 20551 16831 20867 16832
rect 28393 16896 28709 16897
rect 28393 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28639 16896
rect 28703 16832 28709 16896
rect 28393 16831 28709 16832
rect 8788 16352 9104 16353
rect 8788 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8954 16352
rect 9018 16288 9034 16352
rect 9098 16288 9104 16352
rect 8788 16287 9104 16288
rect 16630 16352 16946 16353
rect 16630 16288 16636 16352
rect 16700 16288 16716 16352
rect 16780 16288 16796 16352
rect 16860 16288 16876 16352
rect 16940 16288 16946 16352
rect 16630 16287 16946 16288
rect 24472 16352 24788 16353
rect 24472 16288 24478 16352
rect 24542 16288 24558 16352
rect 24622 16288 24638 16352
rect 24702 16288 24718 16352
rect 24782 16288 24788 16352
rect 24472 16287 24788 16288
rect 32314 16352 32630 16353
rect 32314 16288 32320 16352
rect 32384 16288 32400 16352
rect 32464 16288 32480 16352
rect 32544 16288 32560 16352
rect 32624 16288 32630 16352
rect 32314 16287 32630 16288
rect 4867 15808 5183 15809
rect 4867 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5113 15808
rect 5177 15744 5183 15808
rect 4867 15743 5183 15744
rect 12709 15808 13025 15809
rect 12709 15744 12715 15808
rect 12779 15744 12795 15808
rect 12859 15744 12875 15808
rect 12939 15744 12955 15808
rect 13019 15744 13025 15808
rect 12709 15743 13025 15744
rect 20551 15808 20867 15809
rect 20551 15744 20557 15808
rect 20621 15744 20637 15808
rect 20701 15744 20717 15808
rect 20781 15744 20797 15808
rect 20861 15744 20867 15808
rect 20551 15743 20867 15744
rect 28393 15808 28709 15809
rect 28393 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28639 15808
rect 28703 15744 28709 15808
rect 28393 15743 28709 15744
rect 8788 15264 9104 15265
rect 8788 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8954 15264
rect 9018 15200 9034 15264
rect 9098 15200 9104 15264
rect 8788 15199 9104 15200
rect 16630 15264 16946 15265
rect 16630 15200 16636 15264
rect 16700 15200 16716 15264
rect 16780 15200 16796 15264
rect 16860 15200 16876 15264
rect 16940 15200 16946 15264
rect 16630 15199 16946 15200
rect 24472 15264 24788 15265
rect 24472 15200 24478 15264
rect 24542 15200 24558 15264
rect 24622 15200 24638 15264
rect 24702 15200 24718 15264
rect 24782 15200 24788 15264
rect 24472 15199 24788 15200
rect 32314 15264 32630 15265
rect 32314 15200 32320 15264
rect 32384 15200 32400 15264
rect 32464 15200 32480 15264
rect 32544 15200 32560 15264
rect 32624 15200 32630 15264
rect 32314 15199 32630 15200
rect 4867 14720 5183 14721
rect 4867 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5113 14720
rect 5177 14656 5183 14720
rect 4867 14655 5183 14656
rect 12709 14720 13025 14721
rect 12709 14656 12715 14720
rect 12779 14656 12795 14720
rect 12859 14656 12875 14720
rect 12939 14656 12955 14720
rect 13019 14656 13025 14720
rect 12709 14655 13025 14656
rect 20551 14720 20867 14721
rect 20551 14656 20557 14720
rect 20621 14656 20637 14720
rect 20701 14656 20717 14720
rect 20781 14656 20797 14720
rect 20861 14656 20867 14720
rect 20551 14655 20867 14656
rect 28393 14720 28709 14721
rect 28393 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28639 14720
rect 28703 14656 28709 14720
rect 28393 14655 28709 14656
rect 8788 14176 9104 14177
rect 8788 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8954 14176
rect 9018 14112 9034 14176
rect 9098 14112 9104 14176
rect 8788 14111 9104 14112
rect 16630 14176 16946 14177
rect 16630 14112 16636 14176
rect 16700 14112 16716 14176
rect 16780 14112 16796 14176
rect 16860 14112 16876 14176
rect 16940 14112 16946 14176
rect 16630 14111 16946 14112
rect 24472 14176 24788 14177
rect 24472 14112 24478 14176
rect 24542 14112 24558 14176
rect 24622 14112 24638 14176
rect 24702 14112 24718 14176
rect 24782 14112 24788 14176
rect 24472 14111 24788 14112
rect 32314 14176 32630 14177
rect 32314 14112 32320 14176
rect 32384 14112 32400 14176
rect 32464 14112 32480 14176
rect 32544 14112 32560 14176
rect 32624 14112 32630 14176
rect 32314 14111 32630 14112
rect 4867 13632 5183 13633
rect 4867 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5113 13632
rect 5177 13568 5183 13632
rect 4867 13567 5183 13568
rect 12709 13632 13025 13633
rect 12709 13568 12715 13632
rect 12779 13568 12795 13632
rect 12859 13568 12875 13632
rect 12939 13568 12955 13632
rect 13019 13568 13025 13632
rect 12709 13567 13025 13568
rect 20551 13632 20867 13633
rect 20551 13568 20557 13632
rect 20621 13568 20637 13632
rect 20701 13568 20717 13632
rect 20781 13568 20797 13632
rect 20861 13568 20867 13632
rect 20551 13567 20867 13568
rect 28393 13632 28709 13633
rect 28393 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28639 13632
rect 28703 13568 28709 13632
rect 28393 13567 28709 13568
rect 8788 13088 9104 13089
rect 8788 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8954 13088
rect 9018 13024 9034 13088
rect 9098 13024 9104 13088
rect 8788 13023 9104 13024
rect 16630 13088 16946 13089
rect 16630 13024 16636 13088
rect 16700 13024 16716 13088
rect 16780 13024 16796 13088
rect 16860 13024 16876 13088
rect 16940 13024 16946 13088
rect 16630 13023 16946 13024
rect 24472 13088 24788 13089
rect 24472 13024 24478 13088
rect 24542 13024 24558 13088
rect 24622 13024 24638 13088
rect 24702 13024 24718 13088
rect 24782 13024 24788 13088
rect 24472 13023 24788 13024
rect 32314 13088 32630 13089
rect 32314 13024 32320 13088
rect 32384 13024 32400 13088
rect 32464 13024 32480 13088
rect 32544 13024 32560 13088
rect 32624 13024 32630 13088
rect 32314 13023 32630 13024
rect 4867 12544 5183 12545
rect 4867 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5113 12544
rect 5177 12480 5183 12544
rect 4867 12479 5183 12480
rect 12709 12544 13025 12545
rect 12709 12480 12715 12544
rect 12779 12480 12795 12544
rect 12859 12480 12875 12544
rect 12939 12480 12955 12544
rect 13019 12480 13025 12544
rect 12709 12479 13025 12480
rect 20551 12544 20867 12545
rect 20551 12480 20557 12544
rect 20621 12480 20637 12544
rect 20701 12480 20717 12544
rect 20781 12480 20797 12544
rect 20861 12480 20867 12544
rect 20551 12479 20867 12480
rect 28393 12544 28709 12545
rect 28393 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28639 12544
rect 28703 12480 28709 12544
rect 28393 12479 28709 12480
rect 8788 12000 9104 12001
rect 8788 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8954 12000
rect 9018 11936 9034 12000
rect 9098 11936 9104 12000
rect 8788 11935 9104 11936
rect 16630 12000 16946 12001
rect 16630 11936 16636 12000
rect 16700 11936 16716 12000
rect 16780 11936 16796 12000
rect 16860 11936 16876 12000
rect 16940 11936 16946 12000
rect 16630 11935 16946 11936
rect 24472 12000 24788 12001
rect 24472 11936 24478 12000
rect 24542 11936 24558 12000
rect 24622 11936 24638 12000
rect 24702 11936 24718 12000
rect 24782 11936 24788 12000
rect 24472 11935 24788 11936
rect 32314 12000 32630 12001
rect 32314 11936 32320 12000
rect 32384 11936 32400 12000
rect 32464 11936 32480 12000
rect 32544 11936 32560 12000
rect 32624 11936 32630 12000
rect 32314 11935 32630 11936
rect 4867 11456 5183 11457
rect 4867 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5113 11456
rect 5177 11392 5183 11456
rect 4867 11391 5183 11392
rect 12709 11456 13025 11457
rect 12709 11392 12715 11456
rect 12779 11392 12795 11456
rect 12859 11392 12875 11456
rect 12939 11392 12955 11456
rect 13019 11392 13025 11456
rect 12709 11391 13025 11392
rect 20551 11456 20867 11457
rect 20551 11392 20557 11456
rect 20621 11392 20637 11456
rect 20701 11392 20717 11456
rect 20781 11392 20797 11456
rect 20861 11392 20867 11456
rect 20551 11391 20867 11392
rect 28393 11456 28709 11457
rect 28393 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28639 11456
rect 28703 11392 28709 11456
rect 28393 11391 28709 11392
rect 8788 10912 9104 10913
rect 8788 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8954 10912
rect 9018 10848 9034 10912
rect 9098 10848 9104 10912
rect 8788 10847 9104 10848
rect 16630 10912 16946 10913
rect 16630 10848 16636 10912
rect 16700 10848 16716 10912
rect 16780 10848 16796 10912
rect 16860 10848 16876 10912
rect 16940 10848 16946 10912
rect 16630 10847 16946 10848
rect 24472 10912 24788 10913
rect 24472 10848 24478 10912
rect 24542 10848 24558 10912
rect 24622 10848 24638 10912
rect 24702 10848 24718 10912
rect 24782 10848 24788 10912
rect 24472 10847 24788 10848
rect 32314 10912 32630 10913
rect 32314 10848 32320 10912
rect 32384 10848 32400 10912
rect 32464 10848 32480 10912
rect 32544 10848 32560 10912
rect 32624 10848 32630 10912
rect 32314 10847 32630 10848
rect 4867 10368 5183 10369
rect 4867 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5113 10368
rect 5177 10304 5183 10368
rect 4867 10303 5183 10304
rect 12709 10368 13025 10369
rect 12709 10304 12715 10368
rect 12779 10304 12795 10368
rect 12859 10304 12875 10368
rect 12939 10304 12955 10368
rect 13019 10304 13025 10368
rect 12709 10303 13025 10304
rect 20551 10368 20867 10369
rect 20551 10304 20557 10368
rect 20621 10304 20637 10368
rect 20701 10304 20717 10368
rect 20781 10304 20797 10368
rect 20861 10304 20867 10368
rect 20551 10303 20867 10304
rect 28393 10368 28709 10369
rect 28393 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28639 10368
rect 28703 10304 28709 10368
rect 28393 10303 28709 10304
rect 8788 9824 9104 9825
rect 8788 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8954 9824
rect 9018 9760 9034 9824
rect 9098 9760 9104 9824
rect 8788 9759 9104 9760
rect 16630 9824 16946 9825
rect 16630 9760 16636 9824
rect 16700 9760 16716 9824
rect 16780 9760 16796 9824
rect 16860 9760 16876 9824
rect 16940 9760 16946 9824
rect 16630 9759 16946 9760
rect 24472 9824 24788 9825
rect 24472 9760 24478 9824
rect 24542 9760 24558 9824
rect 24622 9760 24638 9824
rect 24702 9760 24718 9824
rect 24782 9760 24788 9824
rect 24472 9759 24788 9760
rect 32314 9824 32630 9825
rect 32314 9760 32320 9824
rect 32384 9760 32400 9824
rect 32464 9760 32480 9824
rect 32544 9760 32560 9824
rect 32624 9760 32630 9824
rect 32314 9759 32630 9760
rect 4867 9280 5183 9281
rect 4867 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5113 9280
rect 5177 9216 5183 9280
rect 4867 9215 5183 9216
rect 12709 9280 13025 9281
rect 12709 9216 12715 9280
rect 12779 9216 12795 9280
rect 12859 9216 12875 9280
rect 12939 9216 12955 9280
rect 13019 9216 13025 9280
rect 12709 9215 13025 9216
rect 20551 9280 20867 9281
rect 20551 9216 20557 9280
rect 20621 9216 20637 9280
rect 20701 9216 20717 9280
rect 20781 9216 20797 9280
rect 20861 9216 20867 9280
rect 20551 9215 20867 9216
rect 28393 9280 28709 9281
rect 28393 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28639 9280
rect 28703 9216 28709 9280
rect 28393 9215 28709 9216
rect 8788 8736 9104 8737
rect 8788 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8954 8736
rect 9018 8672 9034 8736
rect 9098 8672 9104 8736
rect 8788 8671 9104 8672
rect 16630 8736 16946 8737
rect 16630 8672 16636 8736
rect 16700 8672 16716 8736
rect 16780 8672 16796 8736
rect 16860 8672 16876 8736
rect 16940 8672 16946 8736
rect 16630 8671 16946 8672
rect 24472 8736 24788 8737
rect 24472 8672 24478 8736
rect 24542 8672 24558 8736
rect 24622 8672 24638 8736
rect 24702 8672 24718 8736
rect 24782 8672 24788 8736
rect 24472 8671 24788 8672
rect 32314 8736 32630 8737
rect 32314 8672 32320 8736
rect 32384 8672 32400 8736
rect 32464 8672 32480 8736
rect 32544 8672 32560 8736
rect 32624 8672 32630 8736
rect 32314 8671 32630 8672
rect 4867 8192 5183 8193
rect 4867 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5113 8192
rect 5177 8128 5183 8192
rect 4867 8127 5183 8128
rect 12709 8192 13025 8193
rect 12709 8128 12715 8192
rect 12779 8128 12795 8192
rect 12859 8128 12875 8192
rect 12939 8128 12955 8192
rect 13019 8128 13025 8192
rect 12709 8127 13025 8128
rect 20551 8192 20867 8193
rect 20551 8128 20557 8192
rect 20621 8128 20637 8192
rect 20701 8128 20717 8192
rect 20781 8128 20797 8192
rect 20861 8128 20867 8192
rect 20551 8127 20867 8128
rect 28393 8192 28709 8193
rect 28393 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28639 8192
rect 28703 8128 28709 8192
rect 28393 8127 28709 8128
rect 8788 7648 9104 7649
rect 8788 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8954 7648
rect 9018 7584 9034 7648
rect 9098 7584 9104 7648
rect 8788 7583 9104 7584
rect 16630 7648 16946 7649
rect 16630 7584 16636 7648
rect 16700 7584 16716 7648
rect 16780 7584 16796 7648
rect 16860 7584 16876 7648
rect 16940 7584 16946 7648
rect 16630 7583 16946 7584
rect 24472 7648 24788 7649
rect 24472 7584 24478 7648
rect 24542 7584 24558 7648
rect 24622 7584 24638 7648
rect 24702 7584 24718 7648
rect 24782 7584 24788 7648
rect 24472 7583 24788 7584
rect 32314 7648 32630 7649
rect 32314 7584 32320 7648
rect 32384 7584 32400 7648
rect 32464 7584 32480 7648
rect 32544 7584 32560 7648
rect 32624 7584 32630 7648
rect 32314 7583 32630 7584
rect 4867 7104 5183 7105
rect 4867 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5113 7104
rect 5177 7040 5183 7104
rect 4867 7039 5183 7040
rect 12709 7104 13025 7105
rect 12709 7040 12715 7104
rect 12779 7040 12795 7104
rect 12859 7040 12875 7104
rect 12939 7040 12955 7104
rect 13019 7040 13025 7104
rect 12709 7039 13025 7040
rect 20551 7104 20867 7105
rect 20551 7040 20557 7104
rect 20621 7040 20637 7104
rect 20701 7040 20717 7104
rect 20781 7040 20797 7104
rect 20861 7040 20867 7104
rect 20551 7039 20867 7040
rect 28393 7104 28709 7105
rect 28393 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28639 7104
rect 28703 7040 28709 7104
rect 28393 7039 28709 7040
rect 8788 6560 9104 6561
rect 8788 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8954 6560
rect 9018 6496 9034 6560
rect 9098 6496 9104 6560
rect 8788 6495 9104 6496
rect 16630 6560 16946 6561
rect 16630 6496 16636 6560
rect 16700 6496 16716 6560
rect 16780 6496 16796 6560
rect 16860 6496 16876 6560
rect 16940 6496 16946 6560
rect 16630 6495 16946 6496
rect 24472 6560 24788 6561
rect 24472 6496 24478 6560
rect 24542 6496 24558 6560
rect 24622 6496 24638 6560
rect 24702 6496 24718 6560
rect 24782 6496 24788 6560
rect 24472 6495 24788 6496
rect 32314 6560 32630 6561
rect 32314 6496 32320 6560
rect 32384 6496 32400 6560
rect 32464 6496 32480 6560
rect 32544 6496 32560 6560
rect 32624 6496 32630 6560
rect 32314 6495 32630 6496
rect 4867 6016 5183 6017
rect 4867 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5113 6016
rect 5177 5952 5183 6016
rect 4867 5951 5183 5952
rect 12709 6016 13025 6017
rect 12709 5952 12715 6016
rect 12779 5952 12795 6016
rect 12859 5952 12875 6016
rect 12939 5952 12955 6016
rect 13019 5952 13025 6016
rect 12709 5951 13025 5952
rect 20551 6016 20867 6017
rect 20551 5952 20557 6016
rect 20621 5952 20637 6016
rect 20701 5952 20717 6016
rect 20781 5952 20797 6016
rect 20861 5952 20867 6016
rect 20551 5951 20867 5952
rect 28393 6016 28709 6017
rect 28393 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28639 6016
rect 28703 5952 28709 6016
rect 28393 5951 28709 5952
rect 8788 5472 9104 5473
rect 8788 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8954 5472
rect 9018 5408 9034 5472
rect 9098 5408 9104 5472
rect 8788 5407 9104 5408
rect 16630 5472 16946 5473
rect 16630 5408 16636 5472
rect 16700 5408 16716 5472
rect 16780 5408 16796 5472
rect 16860 5408 16876 5472
rect 16940 5408 16946 5472
rect 16630 5407 16946 5408
rect 24472 5472 24788 5473
rect 24472 5408 24478 5472
rect 24542 5408 24558 5472
rect 24622 5408 24638 5472
rect 24702 5408 24718 5472
rect 24782 5408 24788 5472
rect 24472 5407 24788 5408
rect 32314 5472 32630 5473
rect 32314 5408 32320 5472
rect 32384 5408 32400 5472
rect 32464 5408 32480 5472
rect 32544 5408 32560 5472
rect 32624 5408 32630 5472
rect 32314 5407 32630 5408
rect 4867 4928 5183 4929
rect 4867 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5113 4928
rect 5177 4864 5183 4928
rect 4867 4863 5183 4864
rect 12709 4928 13025 4929
rect 12709 4864 12715 4928
rect 12779 4864 12795 4928
rect 12859 4864 12875 4928
rect 12939 4864 12955 4928
rect 13019 4864 13025 4928
rect 12709 4863 13025 4864
rect 20551 4928 20867 4929
rect 20551 4864 20557 4928
rect 20621 4864 20637 4928
rect 20701 4864 20717 4928
rect 20781 4864 20797 4928
rect 20861 4864 20867 4928
rect 20551 4863 20867 4864
rect 28393 4928 28709 4929
rect 28393 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28639 4928
rect 28703 4864 28709 4928
rect 28393 4863 28709 4864
rect 8788 4384 9104 4385
rect 8788 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8954 4384
rect 9018 4320 9034 4384
rect 9098 4320 9104 4384
rect 8788 4319 9104 4320
rect 16630 4384 16946 4385
rect 16630 4320 16636 4384
rect 16700 4320 16716 4384
rect 16780 4320 16796 4384
rect 16860 4320 16876 4384
rect 16940 4320 16946 4384
rect 16630 4319 16946 4320
rect 24472 4384 24788 4385
rect 24472 4320 24478 4384
rect 24542 4320 24558 4384
rect 24622 4320 24638 4384
rect 24702 4320 24718 4384
rect 24782 4320 24788 4384
rect 24472 4319 24788 4320
rect 32314 4384 32630 4385
rect 32314 4320 32320 4384
rect 32384 4320 32400 4384
rect 32464 4320 32480 4384
rect 32544 4320 32560 4384
rect 32624 4320 32630 4384
rect 32314 4319 32630 4320
rect 4867 3840 5183 3841
rect 4867 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5113 3840
rect 5177 3776 5183 3840
rect 4867 3775 5183 3776
rect 12709 3840 13025 3841
rect 12709 3776 12715 3840
rect 12779 3776 12795 3840
rect 12859 3776 12875 3840
rect 12939 3776 12955 3840
rect 13019 3776 13025 3840
rect 12709 3775 13025 3776
rect 20551 3840 20867 3841
rect 20551 3776 20557 3840
rect 20621 3776 20637 3840
rect 20701 3776 20717 3840
rect 20781 3776 20797 3840
rect 20861 3776 20867 3840
rect 20551 3775 20867 3776
rect 28393 3840 28709 3841
rect 28393 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28639 3840
rect 28703 3776 28709 3840
rect 28393 3775 28709 3776
rect 8788 3296 9104 3297
rect 8788 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8954 3296
rect 9018 3232 9034 3296
rect 9098 3232 9104 3296
rect 8788 3231 9104 3232
rect 16630 3296 16946 3297
rect 16630 3232 16636 3296
rect 16700 3232 16716 3296
rect 16780 3232 16796 3296
rect 16860 3232 16876 3296
rect 16940 3232 16946 3296
rect 16630 3231 16946 3232
rect 24472 3296 24788 3297
rect 24472 3232 24478 3296
rect 24542 3232 24558 3296
rect 24622 3232 24638 3296
rect 24702 3232 24718 3296
rect 24782 3232 24788 3296
rect 24472 3231 24788 3232
rect 32314 3296 32630 3297
rect 32314 3232 32320 3296
rect 32384 3232 32400 3296
rect 32464 3232 32480 3296
rect 32544 3232 32560 3296
rect 32624 3232 32630 3296
rect 32314 3231 32630 3232
rect 4867 2752 5183 2753
rect 4867 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5113 2752
rect 5177 2688 5183 2752
rect 4867 2687 5183 2688
rect 12709 2752 13025 2753
rect 12709 2688 12715 2752
rect 12779 2688 12795 2752
rect 12859 2688 12875 2752
rect 12939 2688 12955 2752
rect 13019 2688 13025 2752
rect 12709 2687 13025 2688
rect 20551 2752 20867 2753
rect 20551 2688 20557 2752
rect 20621 2688 20637 2752
rect 20701 2688 20717 2752
rect 20781 2688 20797 2752
rect 20861 2688 20867 2752
rect 20551 2687 20867 2688
rect 28393 2752 28709 2753
rect 28393 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28639 2752
rect 28703 2688 28709 2752
rect 28393 2687 28709 2688
rect 8788 2208 9104 2209
rect 8788 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8954 2208
rect 9018 2144 9034 2208
rect 9098 2144 9104 2208
rect 8788 2143 9104 2144
rect 16630 2208 16946 2209
rect 16630 2144 16636 2208
rect 16700 2144 16716 2208
rect 16780 2144 16796 2208
rect 16860 2144 16876 2208
rect 16940 2144 16946 2208
rect 16630 2143 16946 2144
rect 24472 2208 24788 2209
rect 24472 2144 24478 2208
rect 24542 2144 24558 2208
rect 24622 2144 24638 2208
rect 24702 2144 24718 2208
rect 24782 2144 24788 2208
rect 24472 2143 24788 2144
rect 32314 2208 32630 2209
rect 32314 2144 32320 2208
rect 32384 2144 32400 2208
rect 32464 2144 32480 2208
rect 32544 2144 32560 2208
rect 32624 2144 32630 2208
rect 32314 2143 32630 2144
rect 4867 1664 5183 1665
rect 4867 1600 4873 1664
rect 4937 1600 4953 1664
rect 5017 1600 5033 1664
rect 5097 1600 5113 1664
rect 5177 1600 5183 1664
rect 4867 1599 5183 1600
rect 12709 1664 13025 1665
rect 12709 1600 12715 1664
rect 12779 1600 12795 1664
rect 12859 1600 12875 1664
rect 12939 1600 12955 1664
rect 13019 1600 13025 1664
rect 12709 1599 13025 1600
rect 20551 1664 20867 1665
rect 20551 1600 20557 1664
rect 20621 1600 20637 1664
rect 20701 1600 20717 1664
rect 20781 1600 20797 1664
rect 20861 1600 20867 1664
rect 20551 1599 20867 1600
rect 28393 1664 28709 1665
rect 28393 1600 28399 1664
rect 28463 1600 28479 1664
rect 28543 1600 28559 1664
rect 28623 1600 28639 1664
rect 28703 1600 28709 1664
rect 28393 1599 28709 1600
rect 8788 1120 9104 1121
rect 8788 1056 8794 1120
rect 8858 1056 8874 1120
rect 8938 1056 8954 1120
rect 9018 1056 9034 1120
rect 9098 1056 9104 1120
rect 8788 1055 9104 1056
rect 16630 1120 16946 1121
rect 16630 1056 16636 1120
rect 16700 1056 16716 1120
rect 16780 1056 16796 1120
rect 16860 1056 16876 1120
rect 16940 1056 16946 1120
rect 16630 1055 16946 1056
rect 24472 1120 24788 1121
rect 24472 1056 24478 1120
rect 24542 1056 24558 1120
rect 24622 1056 24638 1120
rect 24702 1056 24718 1120
rect 24782 1056 24788 1120
rect 24472 1055 24788 1056
rect 32314 1120 32630 1121
rect 32314 1056 32320 1120
rect 32384 1056 32400 1120
rect 32464 1056 32480 1120
rect 32544 1056 32560 1120
rect 32624 1056 32630 1120
rect 32314 1055 32630 1056
rect 260 -2240 1366 -1820
rect 260 -3288 680 -2240
rect 18252 -3288 18956 -3178
rect 260 -3302 18956 -3288
rect 260 -3708 18388 -3302
rect 18252 -3734 18388 -3708
rect 18836 -3734 18956 -3302
rect 18252 -3810 18956 -3734
<< via3 >>
rect 8892 21388 8956 21452
rect 9628 21448 9692 21452
rect 9628 21392 9678 21448
rect 9678 21392 9692 21448
rect 9628 21388 9692 21392
rect 11100 21448 11164 21452
rect 11100 21392 11114 21448
rect 11114 21392 11164 21448
rect 11100 21388 11164 21392
rect 11836 21448 11900 21452
rect 11836 21392 11886 21448
rect 11886 21392 11900 21448
rect 11836 21388 11900 21392
rect 13308 21388 13372 21452
rect 14780 21388 14844 21452
rect 15516 21448 15580 21452
rect 15516 21392 15566 21448
rect 15566 21392 15580 21448
rect 15516 21388 15580 21392
rect 16252 21388 16316 21452
rect 17724 21388 17788 21452
rect 18460 21388 18524 21452
rect 19932 21388 19996 21452
rect 21404 21388 21468 21452
rect 22140 21388 22204 21452
rect 23612 21448 23676 21452
rect 23612 21392 23662 21448
rect 23662 21392 23676 21448
rect 23612 21388 23676 21392
rect 24348 21448 24412 21452
rect 24348 21392 24398 21448
rect 24398 21392 24412 21448
rect 24348 21388 24412 21392
rect 25820 21448 25884 21452
rect 25820 21392 25870 21448
rect 25870 21392 25884 21448
rect 25820 21388 25884 21392
rect 27292 21388 27356 21452
rect 28764 21448 28828 21452
rect 28764 21392 28814 21448
rect 28814 21392 28828 21448
rect 28764 21388 28828 21392
rect 30236 21448 30300 21452
rect 30236 21392 30286 21448
rect 30286 21392 30300 21448
rect 30236 21388 30300 21392
rect 14044 21252 14108 21316
rect 16988 21252 17052 21316
rect 20310 21208 20374 21272
rect 33614 21208 33696 21280
rect 26556 20980 26620 21044
rect 28028 20980 28092 21044
rect 29500 20980 29564 21044
rect 5212 20904 5276 20908
rect 5212 20848 5226 20904
rect 5226 20848 5276 20904
rect 5212 20844 5276 20848
rect 20668 20844 20732 20908
rect 8794 20700 8858 20704
rect 8794 20644 8798 20700
rect 8798 20644 8854 20700
rect 8854 20644 8858 20700
rect 8794 20640 8858 20644
rect 8874 20700 8938 20704
rect 8874 20644 8878 20700
rect 8878 20644 8934 20700
rect 8934 20644 8938 20700
rect 8874 20640 8938 20644
rect 8954 20700 9018 20704
rect 8954 20644 8958 20700
rect 8958 20644 9014 20700
rect 9014 20644 9018 20700
rect 8954 20640 9018 20644
rect 9034 20700 9098 20704
rect 9034 20644 9038 20700
rect 9038 20644 9094 20700
rect 9094 20644 9098 20700
rect 9034 20640 9098 20644
rect 16636 20700 16700 20704
rect 16636 20644 16640 20700
rect 16640 20644 16696 20700
rect 16696 20644 16700 20700
rect 16636 20640 16700 20644
rect 16716 20700 16780 20704
rect 16716 20644 16720 20700
rect 16720 20644 16776 20700
rect 16776 20644 16780 20700
rect 16716 20640 16780 20644
rect 16796 20700 16860 20704
rect 16796 20644 16800 20700
rect 16800 20644 16856 20700
rect 16856 20644 16860 20700
rect 16796 20640 16860 20644
rect 16876 20700 16940 20704
rect 16876 20644 16880 20700
rect 16880 20644 16936 20700
rect 16936 20644 16940 20700
rect 16876 20640 16940 20644
rect 24478 20700 24542 20704
rect 24478 20644 24482 20700
rect 24482 20644 24538 20700
rect 24538 20644 24542 20700
rect 24478 20640 24542 20644
rect 24558 20700 24622 20704
rect 24558 20644 24562 20700
rect 24562 20644 24618 20700
rect 24618 20644 24622 20700
rect 24558 20640 24622 20644
rect 24638 20700 24702 20704
rect 24638 20644 24642 20700
rect 24642 20644 24698 20700
rect 24698 20644 24702 20700
rect 24638 20640 24702 20644
rect 24718 20700 24782 20704
rect 24718 20644 24722 20700
rect 24722 20644 24778 20700
rect 24778 20644 24782 20700
rect 24718 20640 24782 20644
rect 32320 20700 32384 20704
rect 32320 20644 32324 20700
rect 32324 20644 32380 20700
rect 32380 20644 32384 20700
rect 32320 20640 32384 20644
rect 32400 20700 32464 20704
rect 32400 20644 32404 20700
rect 32404 20644 32460 20700
rect 32460 20644 32464 20700
rect 32400 20640 32464 20644
rect 32480 20700 32544 20704
rect 32480 20644 32484 20700
rect 32484 20644 32540 20700
rect 32540 20644 32544 20700
rect 32480 20640 32544 20644
rect 32560 20700 32624 20704
rect 32560 20644 32564 20700
rect 32564 20644 32620 20700
rect 32620 20644 32624 20700
rect 32560 20640 32624 20644
rect 2268 20436 2332 20500
rect 3004 20436 3068 20500
rect 3740 20436 3804 20500
rect 4476 20496 4540 20500
rect 4476 20440 4526 20496
rect 4526 20440 4540 20496
rect 4476 20436 4540 20440
rect 5948 20496 6012 20500
rect 5948 20440 5998 20496
rect 5998 20440 6012 20496
rect 5948 20436 6012 20440
rect 22876 20436 22940 20500
rect 12572 20360 12636 20364
rect 12572 20304 12622 20360
rect 12622 20304 12636 20360
rect 12572 20300 12636 20304
rect 4873 20156 4937 20160
rect 4873 20100 4877 20156
rect 4877 20100 4933 20156
rect 4933 20100 4937 20156
rect 4873 20096 4937 20100
rect 4953 20156 5017 20160
rect 4953 20100 4957 20156
rect 4957 20100 5013 20156
rect 5013 20100 5017 20156
rect 4953 20096 5017 20100
rect 5033 20156 5097 20160
rect 5033 20100 5037 20156
rect 5037 20100 5093 20156
rect 5093 20100 5097 20156
rect 5033 20096 5097 20100
rect 5113 20156 5177 20160
rect 5113 20100 5117 20156
rect 5117 20100 5173 20156
rect 5173 20100 5177 20156
rect 5113 20096 5177 20100
rect 12715 20156 12779 20160
rect 12715 20100 12719 20156
rect 12719 20100 12775 20156
rect 12775 20100 12779 20156
rect 12715 20096 12779 20100
rect 12795 20156 12859 20160
rect 12795 20100 12799 20156
rect 12799 20100 12855 20156
rect 12855 20100 12859 20156
rect 12795 20096 12859 20100
rect 12875 20156 12939 20160
rect 12875 20100 12879 20156
rect 12879 20100 12935 20156
rect 12935 20100 12939 20156
rect 12875 20096 12939 20100
rect 12955 20156 13019 20160
rect 12955 20100 12959 20156
rect 12959 20100 13015 20156
rect 13015 20100 13019 20156
rect 12955 20096 13019 20100
rect 20557 20156 20621 20160
rect 20557 20100 20561 20156
rect 20561 20100 20617 20156
rect 20617 20100 20621 20156
rect 20557 20096 20621 20100
rect 20637 20156 20701 20160
rect 20637 20100 20641 20156
rect 20641 20100 20697 20156
rect 20697 20100 20701 20156
rect 20637 20096 20701 20100
rect 20717 20156 20781 20160
rect 20717 20100 20721 20156
rect 20721 20100 20777 20156
rect 20777 20100 20781 20156
rect 20717 20096 20781 20100
rect 20797 20156 20861 20160
rect 20797 20100 20801 20156
rect 20801 20100 20857 20156
rect 20857 20100 20861 20156
rect 20797 20096 20861 20100
rect 28399 20156 28463 20160
rect 28399 20100 28403 20156
rect 28403 20100 28459 20156
rect 28459 20100 28463 20156
rect 28399 20096 28463 20100
rect 28479 20156 28543 20160
rect 28479 20100 28483 20156
rect 28483 20100 28539 20156
rect 28539 20100 28543 20156
rect 28479 20096 28543 20100
rect 28559 20156 28623 20160
rect 28559 20100 28563 20156
rect 28563 20100 28619 20156
rect 28619 20100 28623 20156
rect 28559 20096 28623 20100
rect 28639 20156 28703 20160
rect 28639 20100 28643 20156
rect 28643 20100 28699 20156
rect 28699 20100 28703 20156
rect 28639 20096 28703 20100
rect 1532 20088 1596 20092
rect 1532 20032 1582 20088
rect 1582 20032 1596 20088
rect 1532 20028 1596 20032
rect 6684 20088 6748 20092
rect 6684 20032 6734 20088
rect 6734 20032 6748 20088
rect 6684 20028 6748 20032
rect 7420 20088 7484 20092
rect 7420 20032 7470 20088
rect 7470 20032 7484 20088
rect 7420 20028 7484 20032
rect 8156 20088 8220 20092
rect 8156 20032 8206 20088
rect 8206 20032 8220 20088
rect 8156 20028 8220 20032
rect 10364 20028 10428 20092
rect 8794 19612 8858 19616
rect 8794 19556 8798 19612
rect 8798 19556 8854 19612
rect 8854 19556 8858 19612
rect 8794 19552 8858 19556
rect 8874 19612 8938 19616
rect 8874 19556 8878 19612
rect 8878 19556 8934 19612
rect 8934 19556 8938 19612
rect 8874 19552 8938 19556
rect 8954 19612 9018 19616
rect 8954 19556 8958 19612
rect 8958 19556 9014 19612
rect 9014 19556 9018 19612
rect 8954 19552 9018 19556
rect 9034 19612 9098 19616
rect 9034 19556 9038 19612
rect 9038 19556 9094 19612
rect 9094 19556 9098 19612
rect 9034 19552 9098 19556
rect 16636 19612 16700 19616
rect 16636 19556 16640 19612
rect 16640 19556 16696 19612
rect 16696 19556 16700 19612
rect 16636 19552 16700 19556
rect 16716 19612 16780 19616
rect 16716 19556 16720 19612
rect 16720 19556 16776 19612
rect 16776 19556 16780 19612
rect 16716 19552 16780 19556
rect 16796 19612 16860 19616
rect 16796 19556 16800 19612
rect 16800 19556 16856 19612
rect 16856 19556 16860 19612
rect 16796 19552 16860 19556
rect 16876 19612 16940 19616
rect 16876 19556 16880 19612
rect 16880 19556 16936 19612
rect 16936 19556 16940 19612
rect 16876 19552 16940 19556
rect 24478 19612 24542 19616
rect 24478 19556 24482 19612
rect 24482 19556 24538 19612
rect 24538 19556 24542 19612
rect 24478 19552 24542 19556
rect 24558 19612 24622 19616
rect 24558 19556 24562 19612
rect 24562 19556 24618 19612
rect 24618 19556 24622 19612
rect 24558 19552 24622 19556
rect 24638 19612 24702 19616
rect 24638 19556 24642 19612
rect 24642 19556 24698 19612
rect 24698 19556 24702 19612
rect 24638 19552 24702 19556
rect 24718 19612 24782 19616
rect 24718 19556 24722 19612
rect 24722 19556 24778 19612
rect 24778 19556 24782 19612
rect 24718 19552 24782 19556
rect 32320 19612 32384 19616
rect 32320 19556 32324 19612
rect 32324 19556 32380 19612
rect 32380 19556 32384 19612
rect 32320 19552 32384 19556
rect 32400 19612 32464 19616
rect 32400 19556 32404 19612
rect 32404 19556 32460 19612
rect 32460 19556 32464 19612
rect 32400 19552 32464 19556
rect 32480 19612 32544 19616
rect 32480 19556 32484 19612
rect 32484 19556 32540 19612
rect 32540 19556 32544 19612
rect 32480 19552 32544 19556
rect 32560 19612 32624 19616
rect 32560 19556 32564 19612
rect 32564 19556 32620 19612
rect 32620 19556 32624 19612
rect 32560 19552 32624 19556
rect 4873 19068 4937 19072
rect 4873 19012 4877 19068
rect 4877 19012 4933 19068
rect 4933 19012 4937 19068
rect 4873 19008 4937 19012
rect 4953 19068 5017 19072
rect 4953 19012 4957 19068
rect 4957 19012 5013 19068
rect 5013 19012 5017 19068
rect 4953 19008 5017 19012
rect 5033 19068 5097 19072
rect 5033 19012 5037 19068
rect 5037 19012 5093 19068
rect 5093 19012 5097 19068
rect 5033 19008 5097 19012
rect 5113 19068 5177 19072
rect 5113 19012 5117 19068
rect 5117 19012 5173 19068
rect 5173 19012 5177 19068
rect 5113 19008 5177 19012
rect 12715 19068 12779 19072
rect 12715 19012 12719 19068
rect 12719 19012 12775 19068
rect 12775 19012 12779 19068
rect 12715 19008 12779 19012
rect 12795 19068 12859 19072
rect 12795 19012 12799 19068
rect 12799 19012 12855 19068
rect 12855 19012 12859 19068
rect 12795 19008 12859 19012
rect 12875 19068 12939 19072
rect 12875 19012 12879 19068
rect 12879 19012 12935 19068
rect 12935 19012 12939 19068
rect 12875 19008 12939 19012
rect 12955 19068 13019 19072
rect 12955 19012 12959 19068
rect 12959 19012 13015 19068
rect 13015 19012 13019 19068
rect 12955 19008 13019 19012
rect 20557 19068 20621 19072
rect 20557 19012 20561 19068
rect 20561 19012 20617 19068
rect 20617 19012 20621 19068
rect 20557 19008 20621 19012
rect 20637 19068 20701 19072
rect 20637 19012 20641 19068
rect 20641 19012 20697 19068
rect 20697 19012 20701 19068
rect 20637 19008 20701 19012
rect 20717 19068 20781 19072
rect 20717 19012 20721 19068
rect 20721 19012 20777 19068
rect 20777 19012 20781 19068
rect 20717 19008 20781 19012
rect 20797 19068 20861 19072
rect 20797 19012 20801 19068
rect 20801 19012 20857 19068
rect 20857 19012 20861 19068
rect 20797 19008 20861 19012
rect 28399 19068 28463 19072
rect 28399 19012 28403 19068
rect 28403 19012 28459 19068
rect 28459 19012 28463 19068
rect 28399 19008 28463 19012
rect 28479 19068 28543 19072
rect 28479 19012 28483 19068
rect 28483 19012 28539 19068
rect 28539 19012 28543 19068
rect 28479 19008 28543 19012
rect 28559 19068 28623 19072
rect 28559 19012 28563 19068
rect 28563 19012 28619 19068
rect 28619 19012 28623 19068
rect 28559 19008 28623 19012
rect 28639 19068 28703 19072
rect 28639 19012 28643 19068
rect 28643 19012 28699 19068
rect 28699 19012 28703 19068
rect 28639 19008 28703 19012
rect 8794 18524 8858 18528
rect 8794 18468 8798 18524
rect 8798 18468 8854 18524
rect 8854 18468 8858 18524
rect 8794 18464 8858 18468
rect 8874 18524 8938 18528
rect 8874 18468 8878 18524
rect 8878 18468 8934 18524
rect 8934 18468 8938 18524
rect 8874 18464 8938 18468
rect 8954 18524 9018 18528
rect 8954 18468 8958 18524
rect 8958 18468 9014 18524
rect 9014 18468 9018 18524
rect 8954 18464 9018 18468
rect 9034 18524 9098 18528
rect 9034 18468 9038 18524
rect 9038 18468 9094 18524
rect 9094 18468 9098 18524
rect 9034 18464 9098 18468
rect 16636 18524 16700 18528
rect 16636 18468 16640 18524
rect 16640 18468 16696 18524
rect 16696 18468 16700 18524
rect 16636 18464 16700 18468
rect 16716 18524 16780 18528
rect 16716 18468 16720 18524
rect 16720 18468 16776 18524
rect 16776 18468 16780 18524
rect 16716 18464 16780 18468
rect 16796 18524 16860 18528
rect 16796 18468 16800 18524
rect 16800 18468 16856 18524
rect 16856 18468 16860 18524
rect 16796 18464 16860 18468
rect 16876 18524 16940 18528
rect 16876 18468 16880 18524
rect 16880 18468 16936 18524
rect 16936 18468 16940 18524
rect 16876 18464 16940 18468
rect 24478 18524 24542 18528
rect 24478 18468 24482 18524
rect 24482 18468 24538 18524
rect 24538 18468 24542 18524
rect 24478 18464 24542 18468
rect 24558 18524 24622 18528
rect 24558 18468 24562 18524
rect 24562 18468 24618 18524
rect 24618 18468 24622 18524
rect 24558 18464 24622 18468
rect 24638 18524 24702 18528
rect 24638 18468 24642 18524
rect 24642 18468 24698 18524
rect 24698 18468 24702 18524
rect 24638 18464 24702 18468
rect 24718 18524 24782 18528
rect 24718 18468 24722 18524
rect 24722 18468 24778 18524
rect 24778 18468 24782 18524
rect 24718 18464 24782 18468
rect 32320 18524 32384 18528
rect 32320 18468 32324 18524
rect 32324 18468 32380 18524
rect 32380 18468 32384 18524
rect 32320 18464 32384 18468
rect 32400 18524 32464 18528
rect 32400 18468 32404 18524
rect 32404 18468 32460 18524
rect 32460 18468 32464 18524
rect 32400 18464 32464 18468
rect 32480 18524 32544 18528
rect 32480 18468 32484 18524
rect 32484 18468 32540 18524
rect 32540 18468 32544 18524
rect 32480 18464 32544 18468
rect 32560 18524 32624 18528
rect 32560 18468 32564 18524
rect 32564 18468 32620 18524
rect 32620 18468 32624 18524
rect 32560 18464 32624 18468
rect 4873 17980 4937 17984
rect 4873 17924 4877 17980
rect 4877 17924 4933 17980
rect 4933 17924 4937 17980
rect 4873 17920 4937 17924
rect 4953 17980 5017 17984
rect 4953 17924 4957 17980
rect 4957 17924 5013 17980
rect 5013 17924 5017 17980
rect 4953 17920 5017 17924
rect 5033 17980 5097 17984
rect 5033 17924 5037 17980
rect 5037 17924 5093 17980
rect 5093 17924 5097 17980
rect 5033 17920 5097 17924
rect 5113 17980 5177 17984
rect 5113 17924 5117 17980
rect 5117 17924 5173 17980
rect 5173 17924 5177 17980
rect 5113 17920 5177 17924
rect 12715 17980 12779 17984
rect 12715 17924 12719 17980
rect 12719 17924 12775 17980
rect 12775 17924 12779 17980
rect 12715 17920 12779 17924
rect 12795 17980 12859 17984
rect 12795 17924 12799 17980
rect 12799 17924 12855 17980
rect 12855 17924 12859 17980
rect 12795 17920 12859 17924
rect 12875 17980 12939 17984
rect 12875 17924 12879 17980
rect 12879 17924 12935 17980
rect 12935 17924 12939 17980
rect 12875 17920 12939 17924
rect 12955 17980 13019 17984
rect 12955 17924 12959 17980
rect 12959 17924 13015 17980
rect 13015 17924 13019 17980
rect 12955 17920 13019 17924
rect 20557 17980 20621 17984
rect 20557 17924 20561 17980
rect 20561 17924 20617 17980
rect 20617 17924 20621 17980
rect 20557 17920 20621 17924
rect 20637 17980 20701 17984
rect 20637 17924 20641 17980
rect 20641 17924 20697 17980
rect 20697 17924 20701 17980
rect 20637 17920 20701 17924
rect 20717 17980 20781 17984
rect 20717 17924 20721 17980
rect 20721 17924 20777 17980
rect 20777 17924 20781 17980
rect 20717 17920 20781 17924
rect 20797 17980 20861 17984
rect 20797 17924 20801 17980
rect 20801 17924 20857 17980
rect 20857 17924 20861 17980
rect 20797 17920 20861 17924
rect 28399 17980 28463 17984
rect 28399 17924 28403 17980
rect 28403 17924 28459 17980
rect 28459 17924 28463 17980
rect 28399 17920 28463 17924
rect 28479 17980 28543 17984
rect 28479 17924 28483 17980
rect 28483 17924 28539 17980
rect 28539 17924 28543 17980
rect 28479 17920 28543 17924
rect 28559 17980 28623 17984
rect 28559 17924 28563 17980
rect 28563 17924 28619 17980
rect 28619 17924 28623 17980
rect 28559 17920 28623 17924
rect 28639 17980 28703 17984
rect 28639 17924 28643 17980
rect 28643 17924 28699 17980
rect 28699 17924 28703 17980
rect 28639 17920 28703 17924
rect 8794 17436 8858 17440
rect 8794 17380 8798 17436
rect 8798 17380 8854 17436
rect 8854 17380 8858 17436
rect 8794 17376 8858 17380
rect 8874 17436 8938 17440
rect 8874 17380 8878 17436
rect 8878 17380 8934 17436
rect 8934 17380 8938 17436
rect 8874 17376 8938 17380
rect 8954 17436 9018 17440
rect 8954 17380 8958 17436
rect 8958 17380 9014 17436
rect 9014 17380 9018 17436
rect 8954 17376 9018 17380
rect 9034 17436 9098 17440
rect 9034 17380 9038 17436
rect 9038 17380 9094 17436
rect 9094 17380 9098 17436
rect 9034 17376 9098 17380
rect 16636 17436 16700 17440
rect 16636 17380 16640 17436
rect 16640 17380 16696 17436
rect 16696 17380 16700 17436
rect 16636 17376 16700 17380
rect 16716 17436 16780 17440
rect 16716 17380 16720 17436
rect 16720 17380 16776 17436
rect 16776 17380 16780 17436
rect 16716 17376 16780 17380
rect 16796 17436 16860 17440
rect 16796 17380 16800 17436
rect 16800 17380 16856 17436
rect 16856 17380 16860 17436
rect 16796 17376 16860 17380
rect 16876 17436 16940 17440
rect 16876 17380 16880 17436
rect 16880 17380 16936 17436
rect 16936 17380 16940 17436
rect 16876 17376 16940 17380
rect 24478 17436 24542 17440
rect 24478 17380 24482 17436
rect 24482 17380 24538 17436
rect 24538 17380 24542 17436
rect 24478 17376 24542 17380
rect 24558 17436 24622 17440
rect 24558 17380 24562 17436
rect 24562 17380 24618 17436
rect 24618 17380 24622 17436
rect 24558 17376 24622 17380
rect 24638 17436 24702 17440
rect 24638 17380 24642 17436
rect 24642 17380 24698 17436
rect 24698 17380 24702 17436
rect 24638 17376 24702 17380
rect 24718 17436 24782 17440
rect 24718 17380 24722 17436
rect 24722 17380 24778 17436
rect 24778 17380 24782 17436
rect 24718 17376 24782 17380
rect 32320 17436 32384 17440
rect 32320 17380 32324 17436
rect 32324 17380 32380 17436
rect 32380 17380 32384 17436
rect 32320 17376 32384 17380
rect 32400 17436 32464 17440
rect 32400 17380 32404 17436
rect 32404 17380 32460 17436
rect 32460 17380 32464 17436
rect 32400 17376 32464 17380
rect 32480 17436 32544 17440
rect 32480 17380 32484 17436
rect 32484 17380 32540 17436
rect 32540 17380 32544 17436
rect 32480 17376 32544 17380
rect 32560 17436 32624 17440
rect 32560 17380 32564 17436
rect 32564 17380 32620 17436
rect 32620 17380 32624 17436
rect 32560 17376 32624 17380
rect 4873 16892 4937 16896
rect 4873 16836 4877 16892
rect 4877 16836 4933 16892
rect 4933 16836 4937 16892
rect 4873 16832 4937 16836
rect 4953 16892 5017 16896
rect 4953 16836 4957 16892
rect 4957 16836 5013 16892
rect 5013 16836 5017 16892
rect 4953 16832 5017 16836
rect 5033 16892 5097 16896
rect 5033 16836 5037 16892
rect 5037 16836 5093 16892
rect 5093 16836 5097 16892
rect 5033 16832 5097 16836
rect 5113 16892 5177 16896
rect 5113 16836 5117 16892
rect 5117 16836 5173 16892
rect 5173 16836 5177 16892
rect 5113 16832 5177 16836
rect 12715 16892 12779 16896
rect 12715 16836 12719 16892
rect 12719 16836 12775 16892
rect 12775 16836 12779 16892
rect 12715 16832 12779 16836
rect 12795 16892 12859 16896
rect 12795 16836 12799 16892
rect 12799 16836 12855 16892
rect 12855 16836 12859 16892
rect 12795 16832 12859 16836
rect 12875 16892 12939 16896
rect 12875 16836 12879 16892
rect 12879 16836 12935 16892
rect 12935 16836 12939 16892
rect 12875 16832 12939 16836
rect 12955 16892 13019 16896
rect 12955 16836 12959 16892
rect 12959 16836 13015 16892
rect 13015 16836 13019 16892
rect 12955 16832 13019 16836
rect 20557 16892 20621 16896
rect 20557 16836 20561 16892
rect 20561 16836 20617 16892
rect 20617 16836 20621 16892
rect 20557 16832 20621 16836
rect 20637 16892 20701 16896
rect 20637 16836 20641 16892
rect 20641 16836 20697 16892
rect 20697 16836 20701 16892
rect 20637 16832 20701 16836
rect 20717 16892 20781 16896
rect 20717 16836 20721 16892
rect 20721 16836 20777 16892
rect 20777 16836 20781 16892
rect 20717 16832 20781 16836
rect 20797 16892 20861 16896
rect 20797 16836 20801 16892
rect 20801 16836 20857 16892
rect 20857 16836 20861 16892
rect 20797 16832 20861 16836
rect 28399 16892 28463 16896
rect 28399 16836 28403 16892
rect 28403 16836 28459 16892
rect 28459 16836 28463 16892
rect 28399 16832 28463 16836
rect 28479 16892 28543 16896
rect 28479 16836 28483 16892
rect 28483 16836 28539 16892
rect 28539 16836 28543 16892
rect 28479 16832 28543 16836
rect 28559 16892 28623 16896
rect 28559 16836 28563 16892
rect 28563 16836 28619 16892
rect 28619 16836 28623 16892
rect 28559 16832 28623 16836
rect 28639 16892 28703 16896
rect 28639 16836 28643 16892
rect 28643 16836 28699 16892
rect 28699 16836 28703 16892
rect 28639 16832 28703 16836
rect 8794 16348 8858 16352
rect 8794 16292 8798 16348
rect 8798 16292 8854 16348
rect 8854 16292 8858 16348
rect 8794 16288 8858 16292
rect 8874 16348 8938 16352
rect 8874 16292 8878 16348
rect 8878 16292 8934 16348
rect 8934 16292 8938 16348
rect 8874 16288 8938 16292
rect 8954 16348 9018 16352
rect 8954 16292 8958 16348
rect 8958 16292 9014 16348
rect 9014 16292 9018 16348
rect 8954 16288 9018 16292
rect 9034 16348 9098 16352
rect 9034 16292 9038 16348
rect 9038 16292 9094 16348
rect 9094 16292 9098 16348
rect 9034 16288 9098 16292
rect 16636 16348 16700 16352
rect 16636 16292 16640 16348
rect 16640 16292 16696 16348
rect 16696 16292 16700 16348
rect 16636 16288 16700 16292
rect 16716 16348 16780 16352
rect 16716 16292 16720 16348
rect 16720 16292 16776 16348
rect 16776 16292 16780 16348
rect 16716 16288 16780 16292
rect 16796 16348 16860 16352
rect 16796 16292 16800 16348
rect 16800 16292 16856 16348
rect 16856 16292 16860 16348
rect 16796 16288 16860 16292
rect 16876 16348 16940 16352
rect 16876 16292 16880 16348
rect 16880 16292 16936 16348
rect 16936 16292 16940 16348
rect 16876 16288 16940 16292
rect 24478 16348 24542 16352
rect 24478 16292 24482 16348
rect 24482 16292 24538 16348
rect 24538 16292 24542 16348
rect 24478 16288 24542 16292
rect 24558 16348 24622 16352
rect 24558 16292 24562 16348
rect 24562 16292 24618 16348
rect 24618 16292 24622 16348
rect 24558 16288 24622 16292
rect 24638 16348 24702 16352
rect 24638 16292 24642 16348
rect 24642 16292 24698 16348
rect 24698 16292 24702 16348
rect 24638 16288 24702 16292
rect 24718 16348 24782 16352
rect 24718 16292 24722 16348
rect 24722 16292 24778 16348
rect 24778 16292 24782 16348
rect 24718 16288 24782 16292
rect 32320 16348 32384 16352
rect 32320 16292 32324 16348
rect 32324 16292 32380 16348
rect 32380 16292 32384 16348
rect 32320 16288 32384 16292
rect 32400 16348 32464 16352
rect 32400 16292 32404 16348
rect 32404 16292 32460 16348
rect 32460 16292 32464 16348
rect 32400 16288 32464 16292
rect 32480 16348 32544 16352
rect 32480 16292 32484 16348
rect 32484 16292 32540 16348
rect 32540 16292 32544 16348
rect 32480 16288 32544 16292
rect 32560 16348 32624 16352
rect 32560 16292 32564 16348
rect 32564 16292 32620 16348
rect 32620 16292 32624 16348
rect 32560 16288 32624 16292
rect 4873 15804 4937 15808
rect 4873 15748 4877 15804
rect 4877 15748 4933 15804
rect 4933 15748 4937 15804
rect 4873 15744 4937 15748
rect 4953 15804 5017 15808
rect 4953 15748 4957 15804
rect 4957 15748 5013 15804
rect 5013 15748 5017 15804
rect 4953 15744 5017 15748
rect 5033 15804 5097 15808
rect 5033 15748 5037 15804
rect 5037 15748 5093 15804
rect 5093 15748 5097 15804
rect 5033 15744 5097 15748
rect 5113 15804 5177 15808
rect 5113 15748 5117 15804
rect 5117 15748 5173 15804
rect 5173 15748 5177 15804
rect 5113 15744 5177 15748
rect 12715 15804 12779 15808
rect 12715 15748 12719 15804
rect 12719 15748 12775 15804
rect 12775 15748 12779 15804
rect 12715 15744 12779 15748
rect 12795 15804 12859 15808
rect 12795 15748 12799 15804
rect 12799 15748 12855 15804
rect 12855 15748 12859 15804
rect 12795 15744 12859 15748
rect 12875 15804 12939 15808
rect 12875 15748 12879 15804
rect 12879 15748 12935 15804
rect 12935 15748 12939 15804
rect 12875 15744 12939 15748
rect 12955 15804 13019 15808
rect 12955 15748 12959 15804
rect 12959 15748 13015 15804
rect 13015 15748 13019 15804
rect 12955 15744 13019 15748
rect 20557 15804 20621 15808
rect 20557 15748 20561 15804
rect 20561 15748 20617 15804
rect 20617 15748 20621 15804
rect 20557 15744 20621 15748
rect 20637 15804 20701 15808
rect 20637 15748 20641 15804
rect 20641 15748 20697 15804
rect 20697 15748 20701 15804
rect 20637 15744 20701 15748
rect 20717 15804 20781 15808
rect 20717 15748 20721 15804
rect 20721 15748 20777 15804
rect 20777 15748 20781 15804
rect 20717 15744 20781 15748
rect 20797 15804 20861 15808
rect 20797 15748 20801 15804
rect 20801 15748 20857 15804
rect 20857 15748 20861 15804
rect 20797 15744 20861 15748
rect 28399 15804 28463 15808
rect 28399 15748 28403 15804
rect 28403 15748 28459 15804
rect 28459 15748 28463 15804
rect 28399 15744 28463 15748
rect 28479 15804 28543 15808
rect 28479 15748 28483 15804
rect 28483 15748 28539 15804
rect 28539 15748 28543 15804
rect 28479 15744 28543 15748
rect 28559 15804 28623 15808
rect 28559 15748 28563 15804
rect 28563 15748 28619 15804
rect 28619 15748 28623 15804
rect 28559 15744 28623 15748
rect 28639 15804 28703 15808
rect 28639 15748 28643 15804
rect 28643 15748 28699 15804
rect 28699 15748 28703 15804
rect 28639 15744 28703 15748
rect 8794 15260 8858 15264
rect 8794 15204 8798 15260
rect 8798 15204 8854 15260
rect 8854 15204 8858 15260
rect 8794 15200 8858 15204
rect 8874 15260 8938 15264
rect 8874 15204 8878 15260
rect 8878 15204 8934 15260
rect 8934 15204 8938 15260
rect 8874 15200 8938 15204
rect 8954 15260 9018 15264
rect 8954 15204 8958 15260
rect 8958 15204 9014 15260
rect 9014 15204 9018 15260
rect 8954 15200 9018 15204
rect 9034 15260 9098 15264
rect 9034 15204 9038 15260
rect 9038 15204 9094 15260
rect 9094 15204 9098 15260
rect 9034 15200 9098 15204
rect 16636 15260 16700 15264
rect 16636 15204 16640 15260
rect 16640 15204 16696 15260
rect 16696 15204 16700 15260
rect 16636 15200 16700 15204
rect 16716 15260 16780 15264
rect 16716 15204 16720 15260
rect 16720 15204 16776 15260
rect 16776 15204 16780 15260
rect 16716 15200 16780 15204
rect 16796 15260 16860 15264
rect 16796 15204 16800 15260
rect 16800 15204 16856 15260
rect 16856 15204 16860 15260
rect 16796 15200 16860 15204
rect 16876 15260 16940 15264
rect 16876 15204 16880 15260
rect 16880 15204 16936 15260
rect 16936 15204 16940 15260
rect 16876 15200 16940 15204
rect 24478 15260 24542 15264
rect 24478 15204 24482 15260
rect 24482 15204 24538 15260
rect 24538 15204 24542 15260
rect 24478 15200 24542 15204
rect 24558 15260 24622 15264
rect 24558 15204 24562 15260
rect 24562 15204 24618 15260
rect 24618 15204 24622 15260
rect 24558 15200 24622 15204
rect 24638 15260 24702 15264
rect 24638 15204 24642 15260
rect 24642 15204 24698 15260
rect 24698 15204 24702 15260
rect 24638 15200 24702 15204
rect 24718 15260 24782 15264
rect 24718 15204 24722 15260
rect 24722 15204 24778 15260
rect 24778 15204 24782 15260
rect 24718 15200 24782 15204
rect 32320 15260 32384 15264
rect 32320 15204 32324 15260
rect 32324 15204 32380 15260
rect 32380 15204 32384 15260
rect 32320 15200 32384 15204
rect 32400 15260 32464 15264
rect 32400 15204 32404 15260
rect 32404 15204 32460 15260
rect 32460 15204 32464 15260
rect 32400 15200 32464 15204
rect 32480 15260 32544 15264
rect 32480 15204 32484 15260
rect 32484 15204 32540 15260
rect 32540 15204 32544 15260
rect 32480 15200 32544 15204
rect 32560 15260 32624 15264
rect 32560 15204 32564 15260
rect 32564 15204 32620 15260
rect 32620 15204 32624 15260
rect 32560 15200 32624 15204
rect 4873 14716 4937 14720
rect 4873 14660 4877 14716
rect 4877 14660 4933 14716
rect 4933 14660 4937 14716
rect 4873 14656 4937 14660
rect 4953 14716 5017 14720
rect 4953 14660 4957 14716
rect 4957 14660 5013 14716
rect 5013 14660 5017 14716
rect 4953 14656 5017 14660
rect 5033 14716 5097 14720
rect 5033 14660 5037 14716
rect 5037 14660 5093 14716
rect 5093 14660 5097 14716
rect 5033 14656 5097 14660
rect 5113 14716 5177 14720
rect 5113 14660 5117 14716
rect 5117 14660 5173 14716
rect 5173 14660 5177 14716
rect 5113 14656 5177 14660
rect 12715 14716 12779 14720
rect 12715 14660 12719 14716
rect 12719 14660 12775 14716
rect 12775 14660 12779 14716
rect 12715 14656 12779 14660
rect 12795 14716 12859 14720
rect 12795 14660 12799 14716
rect 12799 14660 12855 14716
rect 12855 14660 12859 14716
rect 12795 14656 12859 14660
rect 12875 14716 12939 14720
rect 12875 14660 12879 14716
rect 12879 14660 12935 14716
rect 12935 14660 12939 14716
rect 12875 14656 12939 14660
rect 12955 14716 13019 14720
rect 12955 14660 12959 14716
rect 12959 14660 13015 14716
rect 13015 14660 13019 14716
rect 12955 14656 13019 14660
rect 20557 14716 20621 14720
rect 20557 14660 20561 14716
rect 20561 14660 20617 14716
rect 20617 14660 20621 14716
rect 20557 14656 20621 14660
rect 20637 14716 20701 14720
rect 20637 14660 20641 14716
rect 20641 14660 20697 14716
rect 20697 14660 20701 14716
rect 20637 14656 20701 14660
rect 20717 14716 20781 14720
rect 20717 14660 20721 14716
rect 20721 14660 20777 14716
rect 20777 14660 20781 14716
rect 20717 14656 20781 14660
rect 20797 14716 20861 14720
rect 20797 14660 20801 14716
rect 20801 14660 20857 14716
rect 20857 14660 20861 14716
rect 20797 14656 20861 14660
rect 28399 14716 28463 14720
rect 28399 14660 28403 14716
rect 28403 14660 28459 14716
rect 28459 14660 28463 14716
rect 28399 14656 28463 14660
rect 28479 14716 28543 14720
rect 28479 14660 28483 14716
rect 28483 14660 28539 14716
rect 28539 14660 28543 14716
rect 28479 14656 28543 14660
rect 28559 14716 28623 14720
rect 28559 14660 28563 14716
rect 28563 14660 28619 14716
rect 28619 14660 28623 14716
rect 28559 14656 28623 14660
rect 28639 14716 28703 14720
rect 28639 14660 28643 14716
rect 28643 14660 28699 14716
rect 28699 14660 28703 14716
rect 28639 14656 28703 14660
rect 8794 14172 8858 14176
rect 8794 14116 8798 14172
rect 8798 14116 8854 14172
rect 8854 14116 8858 14172
rect 8794 14112 8858 14116
rect 8874 14172 8938 14176
rect 8874 14116 8878 14172
rect 8878 14116 8934 14172
rect 8934 14116 8938 14172
rect 8874 14112 8938 14116
rect 8954 14172 9018 14176
rect 8954 14116 8958 14172
rect 8958 14116 9014 14172
rect 9014 14116 9018 14172
rect 8954 14112 9018 14116
rect 9034 14172 9098 14176
rect 9034 14116 9038 14172
rect 9038 14116 9094 14172
rect 9094 14116 9098 14172
rect 9034 14112 9098 14116
rect 16636 14172 16700 14176
rect 16636 14116 16640 14172
rect 16640 14116 16696 14172
rect 16696 14116 16700 14172
rect 16636 14112 16700 14116
rect 16716 14172 16780 14176
rect 16716 14116 16720 14172
rect 16720 14116 16776 14172
rect 16776 14116 16780 14172
rect 16716 14112 16780 14116
rect 16796 14172 16860 14176
rect 16796 14116 16800 14172
rect 16800 14116 16856 14172
rect 16856 14116 16860 14172
rect 16796 14112 16860 14116
rect 16876 14172 16940 14176
rect 16876 14116 16880 14172
rect 16880 14116 16936 14172
rect 16936 14116 16940 14172
rect 16876 14112 16940 14116
rect 24478 14172 24542 14176
rect 24478 14116 24482 14172
rect 24482 14116 24538 14172
rect 24538 14116 24542 14172
rect 24478 14112 24542 14116
rect 24558 14172 24622 14176
rect 24558 14116 24562 14172
rect 24562 14116 24618 14172
rect 24618 14116 24622 14172
rect 24558 14112 24622 14116
rect 24638 14172 24702 14176
rect 24638 14116 24642 14172
rect 24642 14116 24698 14172
rect 24698 14116 24702 14172
rect 24638 14112 24702 14116
rect 24718 14172 24782 14176
rect 24718 14116 24722 14172
rect 24722 14116 24778 14172
rect 24778 14116 24782 14172
rect 24718 14112 24782 14116
rect 32320 14172 32384 14176
rect 32320 14116 32324 14172
rect 32324 14116 32380 14172
rect 32380 14116 32384 14172
rect 32320 14112 32384 14116
rect 32400 14172 32464 14176
rect 32400 14116 32404 14172
rect 32404 14116 32460 14172
rect 32460 14116 32464 14172
rect 32400 14112 32464 14116
rect 32480 14172 32544 14176
rect 32480 14116 32484 14172
rect 32484 14116 32540 14172
rect 32540 14116 32544 14172
rect 32480 14112 32544 14116
rect 32560 14172 32624 14176
rect 32560 14116 32564 14172
rect 32564 14116 32620 14172
rect 32620 14116 32624 14172
rect 32560 14112 32624 14116
rect 4873 13628 4937 13632
rect 4873 13572 4877 13628
rect 4877 13572 4933 13628
rect 4933 13572 4937 13628
rect 4873 13568 4937 13572
rect 4953 13628 5017 13632
rect 4953 13572 4957 13628
rect 4957 13572 5013 13628
rect 5013 13572 5017 13628
rect 4953 13568 5017 13572
rect 5033 13628 5097 13632
rect 5033 13572 5037 13628
rect 5037 13572 5093 13628
rect 5093 13572 5097 13628
rect 5033 13568 5097 13572
rect 5113 13628 5177 13632
rect 5113 13572 5117 13628
rect 5117 13572 5173 13628
rect 5173 13572 5177 13628
rect 5113 13568 5177 13572
rect 12715 13628 12779 13632
rect 12715 13572 12719 13628
rect 12719 13572 12775 13628
rect 12775 13572 12779 13628
rect 12715 13568 12779 13572
rect 12795 13628 12859 13632
rect 12795 13572 12799 13628
rect 12799 13572 12855 13628
rect 12855 13572 12859 13628
rect 12795 13568 12859 13572
rect 12875 13628 12939 13632
rect 12875 13572 12879 13628
rect 12879 13572 12935 13628
rect 12935 13572 12939 13628
rect 12875 13568 12939 13572
rect 12955 13628 13019 13632
rect 12955 13572 12959 13628
rect 12959 13572 13015 13628
rect 13015 13572 13019 13628
rect 12955 13568 13019 13572
rect 20557 13628 20621 13632
rect 20557 13572 20561 13628
rect 20561 13572 20617 13628
rect 20617 13572 20621 13628
rect 20557 13568 20621 13572
rect 20637 13628 20701 13632
rect 20637 13572 20641 13628
rect 20641 13572 20697 13628
rect 20697 13572 20701 13628
rect 20637 13568 20701 13572
rect 20717 13628 20781 13632
rect 20717 13572 20721 13628
rect 20721 13572 20777 13628
rect 20777 13572 20781 13628
rect 20717 13568 20781 13572
rect 20797 13628 20861 13632
rect 20797 13572 20801 13628
rect 20801 13572 20857 13628
rect 20857 13572 20861 13628
rect 20797 13568 20861 13572
rect 28399 13628 28463 13632
rect 28399 13572 28403 13628
rect 28403 13572 28459 13628
rect 28459 13572 28463 13628
rect 28399 13568 28463 13572
rect 28479 13628 28543 13632
rect 28479 13572 28483 13628
rect 28483 13572 28539 13628
rect 28539 13572 28543 13628
rect 28479 13568 28543 13572
rect 28559 13628 28623 13632
rect 28559 13572 28563 13628
rect 28563 13572 28619 13628
rect 28619 13572 28623 13628
rect 28559 13568 28623 13572
rect 28639 13628 28703 13632
rect 28639 13572 28643 13628
rect 28643 13572 28699 13628
rect 28699 13572 28703 13628
rect 28639 13568 28703 13572
rect 8794 13084 8858 13088
rect 8794 13028 8798 13084
rect 8798 13028 8854 13084
rect 8854 13028 8858 13084
rect 8794 13024 8858 13028
rect 8874 13084 8938 13088
rect 8874 13028 8878 13084
rect 8878 13028 8934 13084
rect 8934 13028 8938 13084
rect 8874 13024 8938 13028
rect 8954 13084 9018 13088
rect 8954 13028 8958 13084
rect 8958 13028 9014 13084
rect 9014 13028 9018 13084
rect 8954 13024 9018 13028
rect 9034 13084 9098 13088
rect 9034 13028 9038 13084
rect 9038 13028 9094 13084
rect 9094 13028 9098 13084
rect 9034 13024 9098 13028
rect 16636 13084 16700 13088
rect 16636 13028 16640 13084
rect 16640 13028 16696 13084
rect 16696 13028 16700 13084
rect 16636 13024 16700 13028
rect 16716 13084 16780 13088
rect 16716 13028 16720 13084
rect 16720 13028 16776 13084
rect 16776 13028 16780 13084
rect 16716 13024 16780 13028
rect 16796 13084 16860 13088
rect 16796 13028 16800 13084
rect 16800 13028 16856 13084
rect 16856 13028 16860 13084
rect 16796 13024 16860 13028
rect 16876 13084 16940 13088
rect 16876 13028 16880 13084
rect 16880 13028 16936 13084
rect 16936 13028 16940 13084
rect 16876 13024 16940 13028
rect 24478 13084 24542 13088
rect 24478 13028 24482 13084
rect 24482 13028 24538 13084
rect 24538 13028 24542 13084
rect 24478 13024 24542 13028
rect 24558 13084 24622 13088
rect 24558 13028 24562 13084
rect 24562 13028 24618 13084
rect 24618 13028 24622 13084
rect 24558 13024 24622 13028
rect 24638 13084 24702 13088
rect 24638 13028 24642 13084
rect 24642 13028 24698 13084
rect 24698 13028 24702 13084
rect 24638 13024 24702 13028
rect 24718 13084 24782 13088
rect 24718 13028 24722 13084
rect 24722 13028 24778 13084
rect 24778 13028 24782 13084
rect 24718 13024 24782 13028
rect 32320 13084 32384 13088
rect 32320 13028 32324 13084
rect 32324 13028 32380 13084
rect 32380 13028 32384 13084
rect 32320 13024 32384 13028
rect 32400 13084 32464 13088
rect 32400 13028 32404 13084
rect 32404 13028 32460 13084
rect 32460 13028 32464 13084
rect 32400 13024 32464 13028
rect 32480 13084 32544 13088
rect 32480 13028 32484 13084
rect 32484 13028 32540 13084
rect 32540 13028 32544 13084
rect 32480 13024 32544 13028
rect 32560 13084 32624 13088
rect 32560 13028 32564 13084
rect 32564 13028 32620 13084
rect 32620 13028 32624 13084
rect 32560 13024 32624 13028
rect 4873 12540 4937 12544
rect 4873 12484 4877 12540
rect 4877 12484 4933 12540
rect 4933 12484 4937 12540
rect 4873 12480 4937 12484
rect 4953 12540 5017 12544
rect 4953 12484 4957 12540
rect 4957 12484 5013 12540
rect 5013 12484 5017 12540
rect 4953 12480 5017 12484
rect 5033 12540 5097 12544
rect 5033 12484 5037 12540
rect 5037 12484 5093 12540
rect 5093 12484 5097 12540
rect 5033 12480 5097 12484
rect 5113 12540 5177 12544
rect 5113 12484 5117 12540
rect 5117 12484 5173 12540
rect 5173 12484 5177 12540
rect 5113 12480 5177 12484
rect 12715 12540 12779 12544
rect 12715 12484 12719 12540
rect 12719 12484 12775 12540
rect 12775 12484 12779 12540
rect 12715 12480 12779 12484
rect 12795 12540 12859 12544
rect 12795 12484 12799 12540
rect 12799 12484 12855 12540
rect 12855 12484 12859 12540
rect 12795 12480 12859 12484
rect 12875 12540 12939 12544
rect 12875 12484 12879 12540
rect 12879 12484 12935 12540
rect 12935 12484 12939 12540
rect 12875 12480 12939 12484
rect 12955 12540 13019 12544
rect 12955 12484 12959 12540
rect 12959 12484 13015 12540
rect 13015 12484 13019 12540
rect 12955 12480 13019 12484
rect 20557 12540 20621 12544
rect 20557 12484 20561 12540
rect 20561 12484 20617 12540
rect 20617 12484 20621 12540
rect 20557 12480 20621 12484
rect 20637 12540 20701 12544
rect 20637 12484 20641 12540
rect 20641 12484 20697 12540
rect 20697 12484 20701 12540
rect 20637 12480 20701 12484
rect 20717 12540 20781 12544
rect 20717 12484 20721 12540
rect 20721 12484 20777 12540
rect 20777 12484 20781 12540
rect 20717 12480 20781 12484
rect 20797 12540 20861 12544
rect 20797 12484 20801 12540
rect 20801 12484 20857 12540
rect 20857 12484 20861 12540
rect 20797 12480 20861 12484
rect 28399 12540 28463 12544
rect 28399 12484 28403 12540
rect 28403 12484 28459 12540
rect 28459 12484 28463 12540
rect 28399 12480 28463 12484
rect 28479 12540 28543 12544
rect 28479 12484 28483 12540
rect 28483 12484 28539 12540
rect 28539 12484 28543 12540
rect 28479 12480 28543 12484
rect 28559 12540 28623 12544
rect 28559 12484 28563 12540
rect 28563 12484 28619 12540
rect 28619 12484 28623 12540
rect 28559 12480 28623 12484
rect 28639 12540 28703 12544
rect 28639 12484 28643 12540
rect 28643 12484 28699 12540
rect 28699 12484 28703 12540
rect 28639 12480 28703 12484
rect 8794 11996 8858 12000
rect 8794 11940 8798 11996
rect 8798 11940 8854 11996
rect 8854 11940 8858 11996
rect 8794 11936 8858 11940
rect 8874 11996 8938 12000
rect 8874 11940 8878 11996
rect 8878 11940 8934 11996
rect 8934 11940 8938 11996
rect 8874 11936 8938 11940
rect 8954 11996 9018 12000
rect 8954 11940 8958 11996
rect 8958 11940 9014 11996
rect 9014 11940 9018 11996
rect 8954 11936 9018 11940
rect 9034 11996 9098 12000
rect 9034 11940 9038 11996
rect 9038 11940 9094 11996
rect 9094 11940 9098 11996
rect 9034 11936 9098 11940
rect 16636 11996 16700 12000
rect 16636 11940 16640 11996
rect 16640 11940 16696 11996
rect 16696 11940 16700 11996
rect 16636 11936 16700 11940
rect 16716 11996 16780 12000
rect 16716 11940 16720 11996
rect 16720 11940 16776 11996
rect 16776 11940 16780 11996
rect 16716 11936 16780 11940
rect 16796 11996 16860 12000
rect 16796 11940 16800 11996
rect 16800 11940 16856 11996
rect 16856 11940 16860 11996
rect 16796 11936 16860 11940
rect 16876 11996 16940 12000
rect 16876 11940 16880 11996
rect 16880 11940 16936 11996
rect 16936 11940 16940 11996
rect 16876 11936 16940 11940
rect 24478 11996 24542 12000
rect 24478 11940 24482 11996
rect 24482 11940 24538 11996
rect 24538 11940 24542 11996
rect 24478 11936 24542 11940
rect 24558 11996 24622 12000
rect 24558 11940 24562 11996
rect 24562 11940 24618 11996
rect 24618 11940 24622 11996
rect 24558 11936 24622 11940
rect 24638 11996 24702 12000
rect 24638 11940 24642 11996
rect 24642 11940 24698 11996
rect 24698 11940 24702 11996
rect 24638 11936 24702 11940
rect 24718 11996 24782 12000
rect 24718 11940 24722 11996
rect 24722 11940 24778 11996
rect 24778 11940 24782 11996
rect 24718 11936 24782 11940
rect 32320 11996 32384 12000
rect 32320 11940 32324 11996
rect 32324 11940 32380 11996
rect 32380 11940 32384 11996
rect 32320 11936 32384 11940
rect 32400 11996 32464 12000
rect 32400 11940 32404 11996
rect 32404 11940 32460 11996
rect 32460 11940 32464 11996
rect 32400 11936 32464 11940
rect 32480 11996 32544 12000
rect 32480 11940 32484 11996
rect 32484 11940 32540 11996
rect 32540 11940 32544 11996
rect 32480 11936 32544 11940
rect 32560 11996 32624 12000
rect 32560 11940 32564 11996
rect 32564 11940 32620 11996
rect 32620 11940 32624 11996
rect 32560 11936 32624 11940
rect 4873 11452 4937 11456
rect 4873 11396 4877 11452
rect 4877 11396 4933 11452
rect 4933 11396 4937 11452
rect 4873 11392 4937 11396
rect 4953 11452 5017 11456
rect 4953 11396 4957 11452
rect 4957 11396 5013 11452
rect 5013 11396 5017 11452
rect 4953 11392 5017 11396
rect 5033 11452 5097 11456
rect 5033 11396 5037 11452
rect 5037 11396 5093 11452
rect 5093 11396 5097 11452
rect 5033 11392 5097 11396
rect 5113 11452 5177 11456
rect 5113 11396 5117 11452
rect 5117 11396 5173 11452
rect 5173 11396 5177 11452
rect 5113 11392 5177 11396
rect 12715 11452 12779 11456
rect 12715 11396 12719 11452
rect 12719 11396 12775 11452
rect 12775 11396 12779 11452
rect 12715 11392 12779 11396
rect 12795 11452 12859 11456
rect 12795 11396 12799 11452
rect 12799 11396 12855 11452
rect 12855 11396 12859 11452
rect 12795 11392 12859 11396
rect 12875 11452 12939 11456
rect 12875 11396 12879 11452
rect 12879 11396 12935 11452
rect 12935 11396 12939 11452
rect 12875 11392 12939 11396
rect 12955 11452 13019 11456
rect 12955 11396 12959 11452
rect 12959 11396 13015 11452
rect 13015 11396 13019 11452
rect 12955 11392 13019 11396
rect 20557 11452 20621 11456
rect 20557 11396 20561 11452
rect 20561 11396 20617 11452
rect 20617 11396 20621 11452
rect 20557 11392 20621 11396
rect 20637 11452 20701 11456
rect 20637 11396 20641 11452
rect 20641 11396 20697 11452
rect 20697 11396 20701 11452
rect 20637 11392 20701 11396
rect 20717 11452 20781 11456
rect 20717 11396 20721 11452
rect 20721 11396 20777 11452
rect 20777 11396 20781 11452
rect 20717 11392 20781 11396
rect 20797 11452 20861 11456
rect 20797 11396 20801 11452
rect 20801 11396 20857 11452
rect 20857 11396 20861 11452
rect 20797 11392 20861 11396
rect 28399 11452 28463 11456
rect 28399 11396 28403 11452
rect 28403 11396 28459 11452
rect 28459 11396 28463 11452
rect 28399 11392 28463 11396
rect 28479 11452 28543 11456
rect 28479 11396 28483 11452
rect 28483 11396 28539 11452
rect 28539 11396 28543 11452
rect 28479 11392 28543 11396
rect 28559 11452 28623 11456
rect 28559 11396 28563 11452
rect 28563 11396 28619 11452
rect 28619 11396 28623 11452
rect 28559 11392 28623 11396
rect 28639 11452 28703 11456
rect 28639 11396 28643 11452
rect 28643 11396 28699 11452
rect 28699 11396 28703 11452
rect 28639 11392 28703 11396
rect 8794 10908 8858 10912
rect 8794 10852 8798 10908
rect 8798 10852 8854 10908
rect 8854 10852 8858 10908
rect 8794 10848 8858 10852
rect 8874 10908 8938 10912
rect 8874 10852 8878 10908
rect 8878 10852 8934 10908
rect 8934 10852 8938 10908
rect 8874 10848 8938 10852
rect 8954 10908 9018 10912
rect 8954 10852 8958 10908
rect 8958 10852 9014 10908
rect 9014 10852 9018 10908
rect 8954 10848 9018 10852
rect 9034 10908 9098 10912
rect 9034 10852 9038 10908
rect 9038 10852 9094 10908
rect 9094 10852 9098 10908
rect 9034 10848 9098 10852
rect 16636 10908 16700 10912
rect 16636 10852 16640 10908
rect 16640 10852 16696 10908
rect 16696 10852 16700 10908
rect 16636 10848 16700 10852
rect 16716 10908 16780 10912
rect 16716 10852 16720 10908
rect 16720 10852 16776 10908
rect 16776 10852 16780 10908
rect 16716 10848 16780 10852
rect 16796 10908 16860 10912
rect 16796 10852 16800 10908
rect 16800 10852 16856 10908
rect 16856 10852 16860 10908
rect 16796 10848 16860 10852
rect 16876 10908 16940 10912
rect 16876 10852 16880 10908
rect 16880 10852 16936 10908
rect 16936 10852 16940 10908
rect 16876 10848 16940 10852
rect 24478 10908 24542 10912
rect 24478 10852 24482 10908
rect 24482 10852 24538 10908
rect 24538 10852 24542 10908
rect 24478 10848 24542 10852
rect 24558 10908 24622 10912
rect 24558 10852 24562 10908
rect 24562 10852 24618 10908
rect 24618 10852 24622 10908
rect 24558 10848 24622 10852
rect 24638 10908 24702 10912
rect 24638 10852 24642 10908
rect 24642 10852 24698 10908
rect 24698 10852 24702 10908
rect 24638 10848 24702 10852
rect 24718 10908 24782 10912
rect 24718 10852 24722 10908
rect 24722 10852 24778 10908
rect 24778 10852 24782 10908
rect 24718 10848 24782 10852
rect 32320 10908 32384 10912
rect 32320 10852 32324 10908
rect 32324 10852 32380 10908
rect 32380 10852 32384 10908
rect 32320 10848 32384 10852
rect 32400 10908 32464 10912
rect 32400 10852 32404 10908
rect 32404 10852 32460 10908
rect 32460 10852 32464 10908
rect 32400 10848 32464 10852
rect 32480 10908 32544 10912
rect 32480 10852 32484 10908
rect 32484 10852 32540 10908
rect 32540 10852 32544 10908
rect 32480 10848 32544 10852
rect 32560 10908 32624 10912
rect 32560 10852 32564 10908
rect 32564 10852 32620 10908
rect 32620 10852 32624 10908
rect 32560 10848 32624 10852
rect 4873 10364 4937 10368
rect 4873 10308 4877 10364
rect 4877 10308 4933 10364
rect 4933 10308 4937 10364
rect 4873 10304 4937 10308
rect 4953 10364 5017 10368
rect 4953 10308 4957 10364
rect 4957 10308 5013 10364
rect 5013 10308 5017 10364
rect 4953 10304 5017 10308
rect 5033 10364 5097 10368
rect 5033 10308 5037 10364
rect 5037 10308 5093 10364
rect 5093 10308 5097 10364
rect 5033 10304 5097 10308
rect 5113 10364 5177 10368
rect 5113 10308 5117 10364
rect 5117 10308 5173 10364
rect 5173 10308 5177 10364
rect 5113 10304 5177 10308
rect 12715 10364 12779 10368
rect 12715 10308 12719 10364
rect 12719 10308 12775 10364
rect 12775 10308 12779 10364
rect 12715 10304 12779 10308
rect 12795 10364 12859 10368
rect 12795 10308 12799 10364
rect 12799 10308 12855 10364
rect 12855 10308 12859 10364
rect 12795 10304 12859 10308
rect 12875 10364 12939 10368
rect 12875 10308 12879 10364
rect 12879 10308 12935 10364
rect 12935 10308 12939 10364
rect 12875 10304 12939 10308
rect 12955 10364 13019 10368
rect 12955 10308 12959 10364
rect 12959 10308 13015 10364
rect 13015 10308 13019 10364
rect 12955 10304 13019 10308
rect 20557 10364 20621 10368
rect 20557 10308 20561 10364
rect 20561 10308 20617 10364
rect 20617 10308 20621 10364
rect 20557 10304 20621 10308
rect 20637 10364 20701 10368
rect 20637 10308 20641 10364
rect 20641 10308 20697 10364
rect 20697 10308 20701 10364
rect 20637 10304 20701 10308
rect 20717 10364 20781 10368
rect 20717 10308 20721 10364
rect 20721 10308 20777 10364
rect 20777 10308 20781 10364
rect 20717 10304 20781 10308
rect 20797 10364 20861 10368
rect 20797 10308 20801 10364
rect 20801 10308 20857 10364
rect 20857 10308 20861 10364
rect 20797 10304 20861 10308
rect 28399 10364 28463 10368
rect 28399 10308 28403 10364
rect 28403 10308 28459 10364
rect 28459 10308 28463 10364
rect 28399 10304 28463 10308
rect 28479 10364 28543 10368
rect 28479 10308 28483 10364
rect 28483 10308 28539 10364
rect 28539 10308 28543 10364
rect 28479 10304 28543 10308
rect 28559 10364 28623 10368
rect 28559 10308 28563 10364
rect 28563 10308 28619 10364
rect 28619 10308 28623 10364
rect 28559 10304 28623 10308
rect 28639 10364 28703 10368
rect 28639 10308 28643 10364
rect 28643 10308 28699 10364
rect 28699 10308 28703 10364
rect 28639 10304 28703 10308
rect 8794 9820 8858 9824
rect 8794 9764 8798 9820
rect 8798 9764 8854 9820
rect 8854 9764 8858 9820
rect 8794 9760 8858 9764
rect 8874 9820 8938 9824
rect 8874 9764 8878 9820
rect 8878 9764 8934 9820
rect 8934 9764 8938 9820
rect 8874 9760 8938 9764
rect 8954 9820 9018 9824
rect 8954 9764 8958 9820
rect 8958 9764 9014 9820
rect 9014 9764 9018 9820
rect 8954 9760 9018 9764
rect 9034 9820 9098 9824
rect 9034 9764 9038 9820
rect 9038 9764 9094 9820
rect 9094 9764 9098 9820
rect 9034 9760 9098 9764
rect 16636 9820 16700 9824
rect 16636 9764 16640 9820
rect 16640 9764 16696 9820
rect 16696 9764 16700 9820
rect 16636 9760 16700 9764
rect 16716 9820 16780 9824
rect 16716 9764 16720 9820
rect 16720 9764 16776 9820
rect 16776 9764 16780 9820
rect 16716 9760 16780 9764
rect 16796 9820 16860 9824
rect 16796 9764 16800 9820
rect 16800 9764 16856 9820
rect 16856 9764 16860 9820
rect 16796 9760 16860 9764
rect 16876 9820 16940 9824
rect 16876 9764 16880 9820
rect 16880 9764 16936 9820
rect 16936 9764 16940 9820
rect 16876 9760 16940 9764
rect 24478 9820 24542 9824
rect 24478 9764 24482 9820
rect 24482 9764 24538 9820
rect 24538 9764 24542 9820
rect 24478 9760 24542 9764
rect 24558 9820 24622 9824
rect 24558 9764 24562 9820
rect 24562 9764 24618 9820
rect 24618 9764 24622 9820
rect 24558 9760 24622 9764
rect 24638 9820 24702 9824
rect 24638 9764 24642 9820
rect 24642 9764 24698 9820
rect 24698 9764 24702 9820
rect 24638 9760 24702 9764
rect 24718 9820 24782 9824
rect 24718 9764 24722 9820
rect 24722 9764 24778 9820
rect 24778 9764 24782 9820
rect 24718 9760 24782 9764
rect 32320 9820 32384 9824
rect 32320 9764 32324 9820
rect 32324 9764 32380 9820
rect 32380 9764 32384 9820
rect 32320 9760 32384 9764
rect 32400 9820 32464 9824
rect 32400 9764 32404 9820
rect 32404 9764 32460 9820
rect 32460 9764 32464 9820
rect 32400 9760 32464 9764
rect 32480 9820 32544 9824
rect 32480 9764 32484 9820
rect 32484 9764 32540 9820
rect 32540 9764 32544 9820
rect 32480 9760 32544 9764
rect 32560 9820 32624 9824
rect 32560 9764 32564 9820
rect 32564 9764 32620 9820
rect 32620 9764 32624 9820
rect 32560 9760 32624 9764
rect 4873 9276 4937 9280
rect 4873 9220 4877 9276
rect 4877 9220 4933 9276
rect 4933 9220 4937 9276
rect 4873 9216 4937 9220
rect 4953 9276 5017 9280
rect 4953 9220 4957 9276
rect 4957 9220 5013 9276
rect 5013 9220 5017 9276
rect 4953 9216 5017 9220
rect 5033 9276 5097 9280
rect 5033 9220 5037 9276
rect 5037 9220 5093 9276
rect 5093 9220 5097 9276
rect 5033 9216 5097 9220
rect 5113 9276 5177 9280
rect 5113 9220 5117 9276
rect 5117 9220 5173 9276
rect 5173 9220 5177 9276
rect 5113 9216 5177 9220
rect 12715 9276 12779 9280
rect 12715 9220 12719 9276
rect 12719 9220 12775 9276
rect 12775 9220 12779 9276
rect 12715 9216 12779 9220
rect 12795 9276 12859 9280
rect 12795 9220 12799 9276
rect 12799 9220 12855 9276
rect 12855 9220 12859 9276
rect 12795 9216 12859 9220
rect 12875 9276 12939 9280
rect 12875 9220 12879 9276
rect 12879 9220 12935 9276
rect 12935 9220 12939 9276
rect 12875 9216 12939 9220
rect 12955 9276 13019 9280
rect 12955 9220 12959 9276
rect 12959 9220 13015 9276
rect 13015 9220 13019 9276
rect 12955 9216 13019 9220
rect 20557 9276 20621 9280
rect 20557 9220 20561 9276
rect 20561 9220 20617 9276
rect 20617 9220 20621 9276
rect 20557 9216 20621 9220
rect 20637 9276 20701 9280
rect 20637 9220 20641 9276
rect 20641 9220 20697 9276
rect 20697 9220 20701 9276
rect 20637 9216 20701 9220
rect 20717 9276 20781 9280
rect 20717 9220 20721 9276
rect 20721 9220 20777 9276
rect 20777 9220 20781 9276
rect 20717 9216 20781 9220
rect 20797 9276 20861 9280
rect 20797 9220 20801 9276
rect 20801 9220 20857 9276
rect 20857 9220 20861 9276
rect 20797 9216 20861 9220
rect 28399 9276 28463 9280
rect 28399 9220 28403 9276
rect 28403 9220 28459 9276
rect 28459 9220 28463 9276
rect 28399 9216 28463 9220
rect 28479 9276 28543 9280
rect 28479 9220 28483 9276
rect 28483 9220 28539 9276
rect 28539 9220 28543 9276
rect 28479 9216 28543 9220
rect 28559 9276 28623 9280
rect 28559 9220 28563 9276
rect 28563 9220 28619 9276
rect 28619 9220 28623 9276
rect 28559 9216 28623 9220
rect 28639 9276 28703 9280
rect 28639 9220 28643 9276
rect 28643 9220 28699 9276
rect 28699 9220 28703 9276
rect 28639 9216 28703 9220
rect 8794 8732 8858 8736
rect 8794 8676 8798 8732
rect 8798 8676 8854 8732
rect 8854 8676 8858 8732
rect 8794 8672 8858 8676
rect 8874 8732 8938 8736
rect 8874 8676 8878 8732
rect 8878 8676 8934 8732
rect 8934 8676 8938 8732
rect 8874 8672 8938 8676
rect 8954 8732 9018 8736
rect 8954 8676 8958 8732
rect 8958 8676 9014 8732
rect 9014 8676 9018 8732
rect 8954 8672 9018 8676
rect 9034 8732 9098 8736
rect 9034 8676 9038 8732
rect 9038 8676 9094 8732
rect 9094 8676 9098 8732
rect 9034 8672 9098 8676
rect 16636 8732 16700 8736
rect 16636 8676 16640 8732
rect 16640 8676 16696 8732
rect 16696 8676 16700 8732
rect 16636 8672 16700 8676
rect 16716 8732 16780 8736
rect 16716 8676 16720 8732
rect 16720 8676 16776 8732
rect 16776 8676 16780 8732
rect 16716 8672 16780 8676
rect 16796 8732 16860 8736
rect 16796 8676 16800 8732
rect 16800 8676 16856 8732
rect 16856 8676 16860 8732
rect 16796 8672 16860 8676
rect 16876 8732 16940 8736
rect 16876 8676 16880 8732
rect 16880 8676 16936 8732
rect 16936 8676 16940 8732
rect 16876 8672 16940 8676
rect 24478 8732 24542 8736
rect 24478 8676 24482 8732
rect 24482 8676 24538 8732
rect 24538 8676 24542 8732
rect 24478 8672 24542 8676
rect 24558 8732 24622 8736
rect 24558 8676 24562 8732
rect 24562 8676 24618 8732
rect 24618 8676 24622 8732
rect 24558 8672 24622 8676
rect 24638 8732 24702 8736
rect 24638 8676 24642 8732
rect 24642 8676 24698 8732
rect 24698 8676 24702 8732
rect 24638 8672 24702 8676
rect 24718 8732 24782 8736
rect 24718 8676 24722 8732
rect 24722 8676 24778 8732
rect 24778 8676 24782 8732
rect 24718 8672 24782 8676
rect 32320 8732 32384 8736
rect 32320 8676 32324 8732
rect 32324 8676 32380 8732
rect 32380 8676 32384 8732
rect 32320 8672 32384 8676
rect 32400 8732 32464 8736
rect 32400 8676 32404 8732
rect 32404 8676 32460 8732
rect 32460 8676 32464 8732
rect 32400 8672 32464 8676
rect 32480 8732 32544 8736
rect 32480 8676 32484 8732
rect 32484 8676 32540 8732
rect 32540 8676 32544 8732
rect 32480 8672 32544 8676
rect 32560 8732 32624 8736
rect 32560 8676 32564 8732
rect 32564 8676 32620 8732
rect 32620 8676 32624 8732
rect 32560 8672 32624 8676
rect 4873 8188 4937 8192
rect 4873 8132 4877 8188
rect 4877 8132 4933 8188
rect 4933 8132 4937 8188
rect 4873 8128 4937 8132
rect 4953 8188 5017 8192
rect 4953 8132 4957 8188
rect 4957 8132 5013 8188
rect 5013 8132 5017 8188
rect 4953 8128 5017 8132
rect 5033 8188 5097 8192
rect 5033 8132 5037 8188
rect 5037 8132 5093 8188
rect 5093 8132 5097 8188
rect 5033 8128 5097 8132
rect 5113 8188 5177 8192
rect 5113 8132 5117 8188
rect 5117 8132 5173 8188
rect 5173 8132 5177 8188
rect 5113 8128 5177 8132
rect 12715 8188 12779 8192
rect 12715 8132 12719 8188
rect 12719 8132 12775 8188
rect 12775 8132 12779 8188
rect 12715 8128 12779 8132
rect 12795 8188 12859 8192
rect 12795 8132 12799 8188
rect 12799 8132 12855 8188
rect 12855 8132 12859 8188
rect 12795 8128 12859 8132
rect 12875 8188 12939 8192
rect 12875 8132 12879 8188
rect 12879 8132 12935 8188
rect 12935 8132 12939 8188
rect 12875 8128 12939 8132
rect 12955 8188 13019 8192
rect 12955 8132 12959 8188
rect 12959 8132 13015 8188
rect 13015 8132 13019 8188
rect 12955 8128 13019 8132
rect 20557 8188 20621 8192
rect 20557 8132 20561 8188
rect 20561 8132 20617 8188
rect 20617 8132 20621 8188
rect 20557 8128 20621 8132
rect 20637 8188 20701 8192
rect 20637 8132 20641 8188
rect 20641 8132 20697 8188
rect 20697 8132 20701 8188
rect 20637 8128 20701 8132
rect 20717 8188 20781 8192
rect 20717 8132 20721 8188
rect 20721 8132 20777 8188
rect 20777 8132 20781 8188
rect 20717 8128 20781 8132
rect 20797 8188 20861 8192
rect 20797 8132 20801 8188
rect 20801 8132 20857 8188
rect 20857 8132 20861 8188
rect 20797 8128 20861 8132
rect 28399 8188 28463 8192
rect 28399 8132 28403 8188
rect 28403 8132 28459 8188
rect 28459 8132 28463 8188
rect 28399 8128 28463 8132
rect 28479 8188 28543 8192
rect 28479 8132 28483 8188
rect 28483 8132 28539 8188
rect 28539 8132 28543 8188
rect 28479 8128 28543 8132
rect 28559 8188 28623 8192
rect 28559 8132 28563 8188
rect 28563 8132 28619 8188
rect 28619 8132 28623 8188
rect 28559 8128 28623 8132
rect 28639 8188 28703 8192
rect 28639 8132 28643 8188
rect 28643 8132 28699 8188
rect 28699 8132 28703 8188
rect 28639 8128 28703 8132
rect 8794 7644 8858 7648
rect 8794 7588 8798 7644
rect 8798 7588 8854 7644
rect 8854 7588 8858 7644
rect 8794 7584 8858 7588
rect 8874 7644 8938 7648
rect 8874 7588 8878 7644
rect 8878 7588 8934 7644
rect 8934 7588 8938 7644
rect 8874 7584 8938 7588
rect 8954 7644 9018 7648
rect 8954 7588 8958 7644
rect 8958 7588 9014 7644
rect 9014 7588 9018 7644
rect 8954 7584 9018 7588
rect 9034 7644 9098 7648
rect 9034 7588 9038 7644
rect 9038 7588 9094 7644
rect 9094 7588 9098 7644
rect 9034 7584 9098 7588
rect 16636 7644 16700 7648
rect 16636 7588 16640 7644
rect 16640 7588 16696 7644
rect 16696 7588 16700 7644
rect 16636 7584 16700 7588
rect 16716 7644 16780 7648
rect 16716 7588 16720 7644
rect 16720 7588 16776 7644
rect 16776 7588 16780 7644
rect 16716 7584 16780 7588
rect 16796 7644 16860 7648
rect 16796 7588 16800 7644
rect 16800 7588 16856 7644
rect 16856 7588 16860 7644
rect 16796 7584 16860 7588
rect 16876 7644 16940 7648
rect 16876 7588 16880 7644
rect 16880 7588 16936 7644
rect 16936 7588 16940 7644
rect 16876 7584 16940 7588
rect 24478 7644 24542 7648
rect 24478 7588 24482 7644
rect 24482 7588 24538 7644
rect 24538 7588 24542 7644
rect 24478 7584 24542 7588
rect 24558 7644 24622 7648
rect 24558 7588 24562 7644
rect 24562 7588 24618 7644
rect 24618 7588 24622 7644
rect 24558 7584 24622 7588
rect 24638 7644 24702 7648
rect 24638 7588 24642 7644
rect 24642 7588 24698 7644
rect 24698 7588 24702 7644
rect 24638 7584 24702 7588
rect 24718 7644 24782 7648
rect 24718 7588 24722 7644
rect 24722 7588 24778 7644
rect 24778 7588 24782 7644
rect 24718 7584 24782 7588
rect 32320 7644 32384 7648
rect 32320 7588 32324 7644
rect 32324 7588 32380 7644
rect 32380 7588 32384 7644
rect 32320 7584 32384 7588
rect 32400 7644 32464 7648
rect 32400 7588 32404 7644
rect 32404 7588 32460 7644
rect 32460 7588 32464 7644
rect 32400 7584 32464 7588
rect 32480 7644 32544 7648
rect 32480 7588 32484 7644
rect 32484 7588 32540 7644
rect 32540 7588 32544 7644
rect 32480 7584 32544 7588
rect 32560 7644 32624 7648
rect 32560 7588 32564 7644
rect 32564 7588 32620 7644
rect 32620 7588 32624 7644
rect 32560 7584 32624 7588
rect 4873 7100 4937 7104
rect 4873 7044 4877 7100
rect 4877 7044 4933 7100
rect 4933 7044 4937 7100
rect 4873 7040 4937 7044
rect 4953 7100 5017 7104
rect 4953 7044 4957 7100
rect 4957 7044 5013 7100
rect 5013 7044 5017 7100
rect 4953 7040 5017 7044
rect 5033 7100 5097 7104
rect 5033 7044 5037 7100
rect 5037 7044 5093 7100
rect 5093 7044 5097 7100
rect 5033 7040 5097 7044
rect 5113 7100 5177 7104
rect 5113 7044 5117 7100
rect 5117 7044 5173 7100
rect 5173 7044 5177 7100
rect 5113 7040 5177 7044
rect 12715 7100 12779 7104
rect 12715 7044 12719 7100
rect 12719 7044 12775 7100
rect 12775 7044 12779 7100
rect 12715 7040 12779 7044
rect 12795 7100 12859 7104
rect 12795 7044 12799 7100
rect 12799 7044 12855 7100
rect 12855 7044 12859 7100
rect 12795 7040 12859 7044
rect 12875 7100 12939 7104
rect 12875 7044 12879 7100
rect 12879 7044 12935 7100
rect 12935 7044 12939 7100
rect 12875 7040 12939 7044
rect 12955 7100 13019 7104
rect 12955 7044 12959 7100
rect 12959 7044 13015 7100
rect 13015 7044 13019 7100
rect 12955 7040 13019 7044
rect 20557 7100 20621 7104
rect 20557 7044 20561 7100
rect 20561 7044 20617 7100
rect 20617 7044 20621 7100
rect 20557 7040 20621 7044
rect 20637 7100 20701 7104
rect 20637 7044 20641 7100
rect 20641 7044 20697 7100
rect 20697 7044 20701 7100
rect 20637 7040 20701 7044
rect 20717 7100 20781 7104
rect 20717 7044 20721 7100
rect 20721 7044 20777 7100
rect 20777 7044 20781 7100
rect 20717 7040 20781 7044
rect 20797 7100 20861 7104
rect 20797 7044 20801 7100
rect 20801 7044 20857 7100
rect 20857 7044 20861 7100
rect 20797 7040 20861 7044
rect 28399 7100 28463 7104
rect 28399 7044 28403 7100
rect 28403 7044 28459 7100
rect 28459 7044 28463 7100
rect 28399 7040 28463 7044
rect 28479 7100 28543 7104
rect 28479 7044 28483 7100
rect 28483 7044 28539 7100
rect 28539 7044 28543 7100
rect 28479 7040 28543 7044
rect 28559 7100 28623 7104
rect 28559 7044 28563 7100
rect 28563 7044 28619 7100
rect 28619 7044 28623 7100
rect 28559 7040 28623 7044
rect 28639 7100 28703 7104
rect 28639 7044 28643 7100
rect 28643 7044 28699 7100
rect 28699 7044 28703 7100
rect 28639 7040 28703 7044
rect 8794 6556 8858 6560
rect 8794 6500 8798 6556
rect 8798 6500 8854 6556
rect 8854 6500 8858 6556
rect 8794 6496 8858 6500
rect 8874 6556 8938 6560
rect 8874 6500 8878 6556
rect 8878 6500 8934 6556
rect 8934 6500 8938 6556
rect 8874 6496 8938 6500
rect 8954 6556 9018 6560
rect 8954 6500 8958 6556
rect 8958 6500 9014 6556
rect 9014 6500 9018 6556
rect 8954 6496 9018 6500
rect 9034 6556 9098 6560
rect 9034 6500 9038 6556
rect 9038 6500 9094 6556
rect 9094 6500 9098 6556
rect 9034 6496 9098 6500
rect 16636 6556 16700 6560
rect 16636 6500 16640 6556
rect 16640 6500 16696 6556
rect 16696 6500 16700 6556
rect 16636 6496 16700 6500
rect 16716 6556 16780 6560
rect 16716 6500 16720 6556
rect 16720 6500 16776 6556
rect 16776 6500 16780 6556
rect 16716 6496 16780 6500
rect 16796 6556 16860 6560
rect 16796 6500 16800 6556
rect 16800 6500 16856 6556
rect 16856 6500 16860 6556
rect 16796 6496 16860 6500
rect 16876 6556 16940 6560
rect 16876 6500 16880 6556
rect 16880 6500 16936 6556
rect 16936 6500 16940 6556
rect 16876 6496 16940 6500
rect 24478 6556 24542 6560
rect 24478 6500 24482 6556
rect 24482 6500 24538 6556
rect 24538 6500 24542 6556
rect 24478 6496 24542 6500
rect 24558 6556 24622 6560
rect 24558 6500 24562 6556
rect 24562 6500 24618 6556
rect 24618 6500 24622 6556
rect 24558 6496 24622 6500
rect 24638 6556 24702 6560
rect 24638 6500 24642 6556
rect 24642 6500 24698 6556
rect 24698 6500 24702 6556
rect 24638 6496 24702 6500
rect 24718 6556 24782 6560
rect 24718 6500 24722 6556
rect 24722 6500 24778 6556
rect 24778 6500 24782 6556
rect 24718 6496 24782 6500
rect 32320 6556 32384 6560
rect 32320 6500 32324 6556
rect 32324 6500 32380 6556
rect 32380 6500 32384 6556
rect 32320 6496 32384 6500
rect 32400 6556 32464 6560
rect 32400 6500 32404 6556
rect 32404 6500 32460 6556
rect 32460 6500 32464 6556
rect 32400 6496 32464 6500
rect 32480 6556 32544 6560
rect 32480 6500 32484 6556
rect 32484 6500 32540 6556
rect 32540 6500 32544 6556
rect 32480 6496 32544 6500
rect 32560 6556 32624 6560
rect 32560 6500 32564 6556
rect 32564 6500 32620 6556
rect 32620 6500 32624 6556
rect 32560 6496 32624 6500
rect 4873 6012 4937 6016
rect 4873 5956 4877 6012
rect 4877 5956 4933 6012
rect 4933 5956 4937 6012
rect 4873 5952 4937 5956
rect 4953 6012 5017 6016
rect 4953 5956 4957 6012
rect 4957 5956 5013 6012
rect 5013 5956 5017 6012
rect 4953 5952 5017 5956
rect 5033 6012 5097 6016
rect 5033 5956 5037 6012
rect 5037 5956 5093 6012
rect 5093 5956 5097 6012
rect 5033 5952 5097 5956
rect 5113 6012 5177 6016
rect 5113 5956 5117 6012
rect 5117 5956 5173 6012
rect 5173 5956 5177 6012
rect 5113 5952 5177 5956
rect 12715 6012 12779 6016
rect 12715 5956 12719 6012
rect 12719 5956 12775 6012
rect 12775 5956 12779 6012
rect 12715 5952 12779 5956
rect 12795 6012 12859 6016
rect 12795 5956 12799 6012
rect 12799 5956 12855 6012
rect 12855 5956 12859 6012
rect 12795 5952 12859 5956
rect 12875 6012 12939 6016
rect 12875 5956 12879 6012
rect 12879 5956 12935 6012
rect 12935 5956 12939 6012
rect 12875 5952 12939 5956
rect 12955 6012 13019 6016
rect 12955 5956 12959 6012
rect 12959 5956 13015 6012
rect 13015 5956 13019 6012
rect 12955 5952 13019 5956
rect 20557 6012 20621 6016
rect 20557 5956 20561 6012
rect 20561 5956 20617 6012
rect 20617 5956 20621 6012
rect 20557 5952 20621 5956
rect 20637 6012 20701 6016
rect 20637 5956 20641 6012
rect 20641 5956 20697 6012
rect 20697 5956 20701 6012
rect 20637 5952 20701 5956
rect 20717 6012 20781 6016
rect 20717 5956 20721 6012
rect 20721 5956 20777 6012
rect 20777 5956 20781 6012
rect 20717 5952 20781 5956
rect 20797 6012 20861 6016
rect 20797 5956 20801 6012
rect 20801 5956 20857 6012
rect 20857 5956 20861 6012
rect 20797 5952 20861 5956
rect 28399 6012 28463 6016
rect 28399 5956 28403 6012
rect 28403 5956 28459 6012
rect 28459 5956 28463 6012
rect 28399 5952 28463 5956
rect 28479 6012 28543 6016
rect 28479 5956 28483 6012
rect 28483 5956 28539 6012
rect 28539 5956 28543 6012
rect 28479 5952 28543 5956
rect 28559 6012 28623 6016
rect 28559 5956 28563 6012
rect 28563 5956 28619 6012
rect 28619 5956 28623 6012
rect 28559 5952 28623 5956
rect 28639 6012 28703 6016
rect 28639 5956 28643 6012
rect 28643 5956 28699 6012
rect 28699 5956 28703 6012
rect 28639 5952 28703 5956
rect 8794 5468 8858 5472
rect 8794 5412 8798 5468
rect 8798 5412 8854 5468
rect 8854 5412 8858 5468
rect 8794 5408 8858 5412
rect 8874 5468 8938 5472
rect 8874 5412 8878 5468
rect 8878 5412 8934 5468
rect 8934 5412 8938 5468
rect 8874 5408 8938 5412
rect 8954 5468 9018 5472
rect 8954 5412 8958 5468
rect 8958 5412 9014 5468
rect 9014 5412 9018 5468
rect 8954 5408 9018 5412
rect 9034 5468 9098 5472
rect 9034 5412 9038 5468
rect 9038 5412 9094 5468
rect 9094 5412 9098 5468
rect 9034 5408 9098 5412
rect 16636 5468 16700 5472
rect 16636 5412 16640 5468
rect 16640 5412 16696 5468
rect 16696 5412 16700 5468
rect 16636 5408 16700 5412
rect 16716 5468 16780 5472
rect 16716 5412 16720 5468
rect 16720 5412 16776 5468
rect 16776 5412 16780 5468
rect 16716 5408 16780 5412
rect 16796 5468 16860 5472
rect 16796 5412 16800 5468
rect 16800 5412 16856 5468
rect 16856 5412 16860 5468
rect 16796 5408 16860 5412
rect 16876 5468 16940 5472
rect 16876 5412 16880 5468
rect 16880 5412 16936 5468
rect 16936 5412 16940 5468
rect 16876 5408 16940 5412
rect 24478 5468 24542 5472
rect 24478 5412 24482 5468
rect 24482 5412 24538 5468
rect 24538 5412 24542 5468
rect 24478 5408 24542 5412
rect 24558 5468 24622 5472
rect 24558 5412 24562 5468
rect 24562 5412 24618 5468
rect 24618 5412 24622 5468
rect 24558 5408 24622 5412
rect 24638 5468 24702 5472
rect 24638 5412 24642 5468
rect 24642 5412 24698 5468
rect 24698 5412 24702 5468
rect 24638 5408 24702 5412
rect 24718 5468 24782 5472
rect 24718 5412 24722 5468
rect 24722 5412 24778 5468
rect 24778 5412 24782 5468
rect 24718 5408 24782 5412
rect 32320 5468 32384 5472
rect 32320 5412 32324 5468
rect 32324 5412 32380 5468
rect 32380 5412 32384 5468
rect 32320 5408 32384 5412
rect 32400 5468 32464 5472
rect 32400 5412 32404 5468
rect 32404 5412 32460 5468
rect 32460 5412 32464 5468
rect 32400 5408 32464 5412
rect 32480 5468 32544 5472
rect 32480 5412 32484 5468
rect 32484 5412 32540 5468
rect 32540 5412 32544 5468
rect 32480 5408 32544 5412
rect 32560 5468 32624 5472
rect 32560 5412 32564 5468
rect 32564 5412 32620 5468
rect 32620 5412 32624 5468
rect 32560 5408 32624 5412
rect 4873 4924 4937 4928
rect 4873 4868 4877 4924
rect 4877 4868 4933 4924
rect 4933 4868 4937 4924
rect 4873 4864 4937 4868
rect 4953 4924 5017 4928
rect 4953 4868 4957 4924
rect 4957 4868 5013 4924
rect 5013 4868 5017 4924
rect 4953 4864 5017 4868
rect 5033 4924 5097 4928
rect 5033 4868 5037 4924
rect 5037 4868 5093 4924
rect 5093 4868 5097 4924
rect 5033 4864 5097 4868
rect 5113 4924 5177 4928
rect 5113 4868 5117 4924
rect 5117 4868 5173 4924
rect 5173 4868 5177 4924
rect 5113 4864 5177 4868
rect 12715 4924 12779 4928
rect 12715 4868 12719 4924
rect 12719 4868 12775 4924
rect 12775 4868 12779 4924
rect 12715 4864 12779 4868
rect 12795 4924 12859 4928
rect 12795 4868 12799 4924
rect 12799 4868 12855 4924
rect 12855 4868 12859 4924
rect 12795 4864 12859 4868
rect 12875 4924 12939 4928
rect 12875 4868 12879 4924
rect 12879 4868 12935 4924
rect 12935 4868 12939 4924
rect 12875 4864 12939 4868
rect 12955 4924 13019 4928
rect 12955 4868 12959 4924
rect 12959 4868 13015 4924
rect 13015 4868 13019 4924
rect 12955 4864 13019 4868
rect 20557 4924 20621 4928
rect 20557 4868 20561 4924
rect 20561 4868 20617 4924
rect 20617 4868 20621 4924
rect 20557 4864 20621 4868
rect 20637 4924 20701 4928
rect 20637 4868 20641 4924
rect 20641 4868 20697 4924
rect 20697 4868 20701 4924
rect 20637 4864 20701 4868
rect 20717 4924 20781 4928
rect 20717 4868 20721 4924
rect 20721 4868 20777 4924
rect 20777 4868 20781 4924
rect 20717 4864 20781 4868
rect 20797 4924 20861 4928
rect 20797 4868 20801 4924
rect 20801 4868 20857 4924
rect 20857 4868 20861 4924
rect 20797 4864 20861 4868
rect 28399 4924 28463 4928
rect 28399 4868 28403 4924
rect 28403 4868 28459 4924
rect 28459 4868 28463 4924
rect 28399 4864 28463 4868
rect 28479 4924 28543 4928
rect 28479 4868 28483 4924
rect 28483 4868 28539 4924
rect 28539 4868 28543 4924
rect 28479 4864 28543 4868
rect 28559 4924 28623 4928
rect 28559 4868 28563 4924
rect 28563 4868 28619 4924
rect 28619 4868 28623 4924
rect 28559 4864 28623 4868
rect 28639 4924 28703 4928
rect 28639 4868 28643 4924
rect 28643 4868 28699 4924
rect 28699 4868 28703 4924
rect 28639 4864 28703 4868
rect 8794 4380 8858 4384
rect 8794 4324 8798 4380
rect 8798 4324 8854 4380
rect 8854 4324 8858 4380
rect 8794 4320 8858 4324
rect 8874 4380 8938 4384
rect 8874 4324 8878 4380
rect 8878 4324 8934 4380
rect 8934 4324 8938 4380
rect 8874 4320 8938 4324
rect 8954 4380 9018 4384
rect 8954 4324 8958 4380
rect 8958 4324 9014 4380
rect 9014 4324 9018 4380
rect 8954 4320 9018 4324
rect 9034 4380 9098 4384
rect 9034 4324 9038 4380
rect 9038 4324 9094 4380
rect 9094 4324 9098 4380
rect 9034 4320 9098 4324
rect 16636 4380 16700 4384
rect 16636 4324 16640 4380
rect 16640 4324 16696 4380
rect 16696 4324 16700 4380
rect 16636 4320 16700 4324
rect 16716 4380 16780 4384
rect 16716 4324 16720 4380
rect 16720 4324 16776 4380
rect 16776 4324 16780 4380
rect 16716 4320 16780 4324
rect 16796 4380 16860 4384
rect 16796 4324 16800 4380
rect 16800 4324 16856 4380
rect 16856 4324 16860 4380
rect 16796 4320 16860 4324
rect 16876 4380 16940 4384
rect 16876 4324 16880 4380
rect 16880 4324 16936 4380
rect 16936 4324 16940 4380
rect 16876 4320 16940 4324
rect 24478 4380 24542 4384
rect 24478 4324 24482 4380
rect 24482 4324 24538 4380
rect 24538 4324 24542 4380
rect 24478 4320 24542 4324
rect 24558 4380 24622 4384
rect 24558 4324 24562 4380
rect 24562 4324 24618 4380
rect 24618 4324 24622 4380
rect 24558 4320 24622 4324
rect 24638 4380 24702 4384
rect 24638 4324 24642 4380
rect 24642 4324 24698 4380
rect 24698 4324 24702 4380
rect 24638 4320 24702 4324
rect 24718 4380 24782 4384
rect 24718 4324 24722 4380
rect 24722 4324 24778 4380
rect 24778 4324 24782 4380
rect 24718 4320 24782 4324
rect 32320 4380 32384 4384
rect 32320 4324 32324 4380
rect 32324 4324 32380 4380
rect 32380 4324 32384 4380
rect 32320 4320 32384 4324
rect 32400 4380 32464 4384
rect 32400 4324 32404 4380
rect 32404 4324 32460 4380
rect 32460 4324 32464 4380
rect 32400 4320 32464 4324
rect 32480 4380 32544 4384
rect 32480 4324 32484 4380
rect 32484 4324 32540 4380
rect 32540 4324 32544 4380
rect 32480 4320 32544 4324
rect 32560 4380 32624 4384
rect 32560 4324 32564 4380
rect 32564 4324 32620 4380
rect 32620 4324 32624 4380
rect 32560 4320 32624 4324
rect 4873 3836 4937 3840
rect 4873 3780 4877 3836
rect 4877 3780 4933 3836
rect 4933 3780 4937 3836
rect 4873 3776 4937 3780
rect 4953 3836 5017 3840
rect 4953 3780 4957 3836
rect 4957 3780 5013 3836
rect 5013 3780 5017 3836
rect 4953 3776 5017 3780
rect 5033 3836 5097 3840
rect 5033 3780 5037 3836
rect 5037 3780 5093 3836
rect 5093 3780 5097 3836
rect 5033 3776 5097 3780
rect 5113 3836 5177 3840
rect 5113 3780 5117 3836
rect 5117 3780 5173 3836
rect 5173 3780 5177 3836
rect 5113 3776 5177 3780
rect 12715 3836 12779 3840
rect 12715 3780 12719 3836
rect 12719 3780 12775 3836
rect 12775 3780 12779 3836
rect 12715 3776 12779 3780
rect 12795 3836 12859 3840
rect 12795 3780 12799 3836
rect 12799 3780 12855 3836
rect 12855 3780 12859 3836
rect 12795 3776 12859 3780
rect 12875 3836 12939 3840
rect 12875 3780 12879 3836
rect 12879 3780 12935 3836
rect 12935 3780 12939 3836
rect 12875 3776 12939 3780
rect 12955 3836 13019 3840
rect 12955 3780 12959 3836
rect 12959 3780 13015 3836
rect 13015 3780 13019 3836
rect 12955 3776 13019 3780
rect 20557 3836 20621 3840
rect 20557 3780 20561 3836
rect 20561 3780 20617 3836
rect 20617 3780 20621 3836
rect 20557 3776 20621 3780
rect 20637 3836 20701 3840
rect 20637 3780 20641 3836
rect 20641 3780 20697 3836
rect 20697 3780 20701 3836
rect 20637 3776 20701 3780
rect 20717 3836 20781 3840
rect 20717 3780 20721 3836
rect 20721 3780 20777 3836
rect 20777 3780 20781 3836
rect 20717 3776 20781 3780
rect 20797 3836 20861 3840
rect 20797 3780 20801 3836
rect 20801 3780 20857 3836
rect 20857 3780 20861 3836
rect 20797 3776 20861 3780
rect 28399 3836 28463 3840
rect 28399 3780 28403 3836
rect 28403 3780 28459 3836
rect 28459 3780 28463 3836
rect 28399 3776 28463 3780
rect 28479 3836 28543 3840
rect 28479 3780 28483 3836
rect 28483 3780 28539 3836
rect 28539 3780 28543 3836
rect 28479 3776 28543 3780
rect 28559 3836 28623 3840
rect 28559 3780 28563 3836
rect 28563 3780 28619 3836
rect 28619 3780 28623 3836
rect 28559 3776 28623 3780
rect 28639 3836 28703 3840
rect 28639 3780 28643 3836
rect 28643 3780 28699 3836
rect 28699 3780 28703 3836
rect 28639 3776 28703 3780
rect 8794 3292 8858 3296
rect 8794 3236 8798 3292
rect 8798 3236 8854 3292
rect 8854 3236 8858 3292
rect 8794 3232 8858 3236
rect 8874 3292 8938 3296
rect 8874 3236 8878 3292
rect 8878 3236 8934 3292
rect 8934 3236 8938 3292
rect 8874 3232 8938 3236
rect 8954 3292 9018 3296
rect 8954 3236 8958 3292
rect 8958 3236 9014 3292
rect 9014 3236 9018 3292
rect 8954 3232 9018 3236
rect 9034 3292 9098 3296
rect 9034 3236 9038 3292
rect 9038 3236 9094 3292
rect 9094 3236 9098 3292
rect 9034 3232 9098 3236
rect 16636 3292 16700 3296
rect 16636 3236 16640 3292
rect 16640 3236 16696 3292
rect 16696 3236 16700 3292
rect 16636 3232 16700 3236
rect 16716 3292 16780 3296
rect 16716 3236 16720 3292
rect 16720 3236 16776 3292
rect 16776 3236 16780 3292
rect 16716 3232 16780 3236
rect 16796 3292 16860 3296
rect 16796 3236 16800 3292
rect 16800 3236 16856 3292
rect 16856 3236 16860 3292
rect 16796 3232 16860 3236
rect 16876 3292 16940 3296
rect 16876 3236 16880 3292
rect 16880 3236 16936 3292
rect 16936 3236 16940 3292
rect 16876 3232 16940 3236
rect 24478 3292 24542 3296
rect 24478 3236 24482 3292
rect 24482 3236 24538 3292
rect 24538 3236 24542 3292
rect 24478 3232 24542 3236
rect 24558 3292 24622 3296
rect 24558 3236 24562 3292
rect 24562 3236 24618 3292
rect 24618 3236 24622 3292
rect 24558 3232 24622 3236
rect 24638 3292 24702 3296
rect 24638 3236 24642 3292
rect 24642 3236 24698 3292
rect 24698 3236 24702 3292
rect 24638 3232 24702 3236
rect 24718 3292 24782 3296
rect 24718 3236 24722 3292
rect 24722 3236 24778 3292
rect 24778 3236 24782 3292
rect 24718 3232 24782 3236
rect 32320 3292 32384 3296
rect 32320 3236 32324 3292
rect 32324 3236 32380 3292
rect 32380 3236 32384 3292
rect 32320 3232 32384 3236
rect 32400 3292 32464 3296
rect 32400 3236 32404 3292
rect 32404 3236 32460 3292
rect 32460 3236 32464 3292
rect 32400 3232 32464 3236
rect 32480 3292 32544 3296
rect 32480 3236 32484 3292
rect 32484 3236 32540 3292
rect 32540 3236 32544 3292
rect 32480 3232 32544 3236
rect 32560 3292 32624 3296
rect 32560 3236 32564 3292
rect 32564 3236 32620 3292
rect 32620 3236 32624 3292
rect 32560 3232 32624 3236
rect 4873 2748 4937 2752
rect 4873 2692 4877 2748
rect 4877 2692 4933 2748
rect 4933 2692 4937 2748
rect 4873 2688 4937 2692
rect 4953 2748 5017 2752
rect 4953 2692 4957 2748
rect 4957 2692 5013 2748
rect 5013 2692 5017 2748
rect 4953 2688 5017 2692
rect 5033 2748 5097 2752
rect 5033 2692 5037 2748
rect 5037 2692 5093 2748
rect 5093 2692 5097 2748
rect 5033 2688 5097 2692
rect 5113 2748 5177 2752
rect 5113 2692 5117 2748
rect 5117 2692 5173 2748
rect 5173 2692 5177 2748
rect 5113 2688 5177 2692
rect 12715 2748 12779 2752
rect 12715 2692 12719 2748
rect 12719 2692 12775 2748
rect 12775 2692 12779 2748
rect 12715 2688 12779 2692
rect 12795 2748 12859 2752
rect 12795 2692 12799 2748
rect 12799 2692 12855 2748
rect 12855 2692 12859 2748
rect 12795 2688 12859 2692
rect 12875 2748 12939 2752
rect 12875 2692 12879 2748
rect 12879 2692 12935 2748
rect 12935 2692 12939 2748
rect 12875 2688 12939 2692
rect 12955 2748 13019 2752
rect 12955 2692 12959 2748
rect 12959 2692 13015 2748
rect 13015 2692 13019 2748
rect 12955 2688 13019 2692
rect 20557 2748 20621 2752
rect 20557 2692 20561 2748
rect 20561 2692 20617 2748
rect 20617 2692 20621 2748
rect 20557 2688 20621 2692
rect 20637 2748 20701 2752
rect 20637 2692 20641 2748
rect 20641 2692 20697 2748
rect 20697 2692 20701 2748
rect 20637 2688 20701 2692
rect 20717 2748 20781 2752
rect 20717 2692 20721 2748
rect 20721 2692 20777 2748
rect 20777 2692 20781 2748
rect 20717 2688 20781 2692
rect 20797 2748 20861 2752
rect 20797 2692 20801 2748
rect 20801 2692 20857 2748
rect 20857 2692 20861 2748
rect 20797 2688 20861 2692
rect 28399 2748 28463 2752
rect 28399 2692 28403 2748
rect 28403 2692 28459 2748
rect 28459 2692 28463 2748
rect 28399 2688 28463 2692
rect 28479 2748 28543 2752
rect 28479 2692 28483 2748
rect 28483 2692 28539 2748
rect 28539 2692 28543 2748
rect 28479 2688 28543 2692
rect 28559 2748 28623 2752
rect 28559 2692 28563 2748
rect 28563 2692 28619 2748
rect 28619 2692 28623 2748
rect 28559 2688 28623 2692
rect 28639 2748 28703 2752
rect 28639 2692 28643 2748
rect 28643 2692 28699 2748
rect 28699 2692 28703 2748
rect 28639 2688 28703 2692
rect 8794 2204 8858 2208
rect 8794 2148 8798 2204
rect 8798 2148 8854 2204
rect 8854 2148 8858 2204
rect 8794 2144 8858 2148
rect 8874 2204 8938 2208
rect 8874 2148 8878 2204
rect 8878 2148 8934 2204
rect 8934 2148 8938 2204
rect 8874 2144 8938 2148
rect 8954 2204 9018 2208
rect 8954 2148 8958 2204
rect 8958 2148 9014 2204
rect 9014 2148 9018 2204
rect 8954 2144 9018 2148
rect 9034 2204 9098 2208
rect 9034 2148 9038 2204
rect 9038 2148 9094 2204
rect 9094 2148 9098 2204
rect 9034 2144 9098 2148
rect 16636 2204 16700 2208
rect 16636 2148 16640 2204
rect 16640 2148 16696 2204
rect 16696 2148 16700 2204
rect 16636 2144 16700 2148
rect 16716 2204 16780 2208
rect 16716 2148 16720 2204
rect 16720 2148 16776 2204
rect 16776 2148 16780 2204
rect 16716 2144 16780 2148
rect 16796 2204 16860 2208
rect 16796 2148 16800 2204
rect 16800 2148 16856 2204
rect 16856 2148 16860 2204
rect 16796 2144 16860 2148
rect 16876 2204 16940 2208
rect 16876 2148 16880 2204
rect 16880 2148 16936 2204
rect 16936 2148 16940 2204
rect 16876 2144 16940 2148
rect 24478 2204 24542 2208
rect 24478 2148 24482 2204
rect 24482 2148 24538 2204
rect 24538 2148 24542 2204
rect 24478 2144 24542 2148
rect 24558 2204 24622 2208
rect 24558 2148 24562 2204
rect 24562 2148 24618 2204
rect 24618 2148 24622 2204
rect 24558 2144 24622 2148
rect 24638 2204 24702 2208
rect 24638 2148 24642 2204
rect 24642 2148 24698 2204
rect 24698 2148 24702 2204
rect 24638 2144 24702 2148
rect 24718 2204 24782 2208
rect 24718 2148 24722 2204
rect 24722 2148 24778 2204
rect 24778 2148 24782 2204
rect 24718 2144 24782 2148
rect 32320 2204 32384 2208
rect 32320 2148 32324 2204
rect 32324 2148 32380 2204
rect 32380 2148 32384 2204
rect 32320 2144 32384 2148
rect 32400 2204 32464 2208
rect 32400 2148 32404 2204
rect 32404 2148 32460 2204
rect 32460 2148 32464 2204
rect 32400 2144 32464 2148
rect 32480 2204 32544 2208
rect 32480 2148 32484 2204
rect 32484 2148 32540 2204
rect 32540 2148 32544 2204
rect 32480 2144 32544 2148
rect 32560 2204 32624 2208
rect 32560 2148 32564 2204
rect 32564 2148 32620 2204
rect 32620 2148 32624 2204
rect 32560 2144 32624 2148
rect 4873 1660 4937 1664
rect 4873 1604 4877 1660
rect 4877 1604 4933 1660
rect 4933 1604 4937 1660
rect 4873 1600 4937 1604
rect 4953 1660 5017 1664
rect 4953 1604 4957 1660
rect 4957 1604 5013 1660
rect 5013 1604 5017 1660
rect 4953 1600 5017 1604
rect 5033 1660 5097 1664
rect 5033 1604 5037 1660
rect 5037 1604 5093 1660
rect 5093 1604 5097 1660
rect 5033 1600 5097 1604
rect 5113 1660 5177 1664
rect 5113 1604 5117 1660
rect 5117 1604 5173 1660
rect 5173 1604 5177 1660
rect 5113 1600 5177 1604
rect 12715 1660 12779 1664
rect 12715 1604 12719 1660
rect 12719 1604 12775 1660
rect 12775 1604 12779 1660
rect 12715 1600 12779 1604
rect 12795 1660 12859 1664
rect 12795 1604 12799 1660
rect 12799 1604 12855 1660
rect 12855 1604 12859 1660
rect 12795 1600 12859 1604
rect 12875 1660 12939 1664
rect 12875 1604 12879 1660
rect 12879 1604 12935 1660
rect 12935 1604 12939 1660
rect 12875 1600 12939 1604
rect 12955 1660 13019 1664
rect 12955 1604 12959 1660
rect 12959 1604 13015 1660
rect 13015 1604 13019 1660
rect 12955 1600 13019 1604
rect 20557 1660 20621 1664
rect 20557 1604 20561 1660
rect 20561 1604 20617 1660
rect 20617 1604 20621 1660
rect 20557 1600 20621 1604
rect 20637 1660 20701 1664
rect 20637 1604 20641 1660
rect 20641 1604 20697 1660
rect 20697 1604 20701 1660
rect 20637 1600 20701 1604
rect 20717 1660 20781 1664
rect 20717 1604 20721 1660
rect 20721 1604 20777 1660
rect 20777 1604 20781 1660
rect 20717 1600 20781 1604
rect 20797 1660 20861 1664
rect 20797 1604 20801 1660
rect 20801 1604 20857 1660
rect 20857 1604 20861 1660
rect 20797 1600 20861 1604
rect 28399 1660 28463 1664
rect 28399 1604 28403 1660
rect 28403 1604 28459 1660
rect 28459 1604 28463 1660
rect 28399 1600 28463 1604
rect 28479 1660 28543 1664
rect 28479 1604 28483 1660
rect 28483 1604 28539 1660
rect 28539 1604 28543 1660
rect 28479 1600 28543 1604
rect 28559 1660 28623 1664
rect 28559 1604 28563 1660
rect 28563 1604 28619 1660
rect 28619 1604 28623 1660
rect 28559 1600 28623 1604
rect 28639 1660 28703 1664
rect 28639 1604 28643 1660
rect 28643 1604 28699 1660
rect 28699 1604 28703 1660
rect 28639 1600 28703 1604
rect 8794 1116 8858 1120
rect 8794 1060 8798 1116
rect 8798 1060 8854 1116
rect 8854 1060 8858 1116
rect 8794 1056 8858 1060
rect 8874 1116 8938 1120
rect 8874 1060 8878 1116
rect 8878 1060 8934 1116
rect 8934 1060 8938 1116
rect 8874 1056 8938 1060
rect 8954 1116 9018 1120
rect 8954 1060 8958 1116
rect 8958 1060 9014 1116
rect 9014 1060 9018 1116
rect 8954 1056 9018 1060
rect 9034 1116 9098 1120
rect 9034 1060 9038 1116
rect 9038 1060 9094 1116
rect 9094 1060 9098 1116
rect 9034 1056 9098 1060
rect 16636 1116 16700 1120
rect 16636 1060 16640 1116
rect 16640 1060 16696 1116
rect 16696 1060 16700 1116
rect 16636 1056 16700 1060
rect 16716 1116 16780 1120
rect 16716 1060 16720 1116
rect 16720 1060 16776 1116
rect 16776 1060 16780 1116
rect 16716 1056 16780 1060
rect 16796 1116 16860 1120
rect 16796 1060 16800 1116
rect 16800 1060 16856 1116
rect 16856 1060 16860 1116
rect 16796 1056 16860 1060
rect 16876 1116 16940 1120
rect 16876 1060 16880 1116
rect 16880 1060 16936 1116
rect 16936 1060 16940 1116
rect 16876 1056 16940 1060
rect 24478 1116 24542 1120
rect 24478 1060 24482 1116
rect 24482 1060 24538 1116
rect 24538 1060 24542 1116
rect 24478 1056 24542 1060
rect 24558 1116 24622 1120
rect 24558 1060 24562 1116
rect 24562 1060 24618 1116
rect 24618 1060 24622 1116
rect 24558 1056 24622 1060
rect 24638 1116 24702 1120
rect 24638 1060 24642 1116
rect 24642 1060 24698 1116
rect 24698 1060 24702 1116
rect 24638 1056 24702 1060
rect 24718 1116 24782 1120
rect 24718 1060 24722 1116
rect 24722 1060 24778 1116
rect 24778 1060 24782 1116
rect 24718 1056 24782 1060
rect 32320 1116 32384 1120
rect 32320 1060 32324 1116
rect 32324 1060 32380 1116
rect 32380 1060 32384 1116
rect 32320 1056 32384 1060
rect 32400 1116 32464 1120
rect 32400 1060 32404 1116
rect 32404 1060 32460 1116
rect 32460 1060 32464 1116
rect 32400 1056 32464 1060
rect 32480 1116 32544 1120
rect 32480 1060 32484 1116
rect 32484 1060 32540 1116
rect 32540 1060 32544 1116
rect 32480 1056 32544 1060
rect 32560 1116 32624 1120
rect 32560 1060 32564 1116
rect 32564 1060 32620 1116
rect 32620 1060 32624 1116
rect 32560 1056 32624 1060
rect 2172 -882 13766 -634
rect 1262 -2636 1526 -2470
rect 2134 -2598 13776 -2342
rect 18388 -3734 18836 -3302
<< metal4 >>
rect 242 20568 562 20626
rect -54 320 590 20568
rect 1534 20093 1594 21760
rect 2270 20501 2330 21760
rect 3006 20501 3066 21760
rect 3742 20501 3802 21760
rect 4478 20501 4538 21760
rect 5214 20909 5274 21760
rect 5211 20908 5277 20909
rect 5211 20844 5212 20908
rect 5276 20844 5277 20908
rect 5211 20843 5277 20844
rect 2267 20500 2333 20501
rect 2267 20436 2268 20500
rect 2332 20436 2333 20500
rect 2267 20435 2333 20436
rect 3003 20500 3069 20501
rect 3003 20436 3004 20500
rect 3068 20436 3069 20500
rect 3003 20435 3069 20436
rect 3739 20500 3805 20501
rect 3739 20436 3740 20500
rect 3804 20436 3805 20500
rect 3739 20435 3805 20436
rect 4475 20500 4541 20501
rect 4475 20436 4476 20500
rect 4540 20436 4541 20500
rect 4475 20435 4541 20436
rect 4865 20160 5185 20720
rect 5950 20501 6010 21760
rect 5947 20500 6013 20501
rect 5947 20436 5948 20500
rect 6012 20436 6013 20500
rect 5947 20435 6013 20436
rect 4865 20096 4873 20160
rect 4937 20096 4953 20160
rect 5017 20096 5033 20160
rect 5097 20096 5113 20160
rect 5177 20096 5185 20160
rect 1531 20092 1597 20093
rect 1531 20028 1532 20092
rect 1596 20028 1597 20092
rect 1531 20027 1597 20028
rect 4865 19072 5185 20096
rect 6686 20093 6746 21760
rect 7422 20093 7482 21760
rect 8158 20093 8218 21760
rect 8894 21453 8954 21760
rect 9630 21453 9690 21760
rect 8891 21452 8957 21453
rect 8891 21388 8892 21452
rect 8956 21388 8957 21452
rect 8891 21387 8957 21388
rect 9627 21452 9693 21453
rect 9627 21388 9628 21452
rect 9692 21388 9693 21452
rect 9627 21387 9693 21388
rect 8786 20704 9106 20720
rect 8786 20640 8794 20704
rect 8858 20640 8874 20704
rect 8938 20640 8954 20704
rect 9018 20640 9034 20704
rect 9098 20640 9106 20704
rect 6683 20092 6749 20093
rect 6683 20028 6684 20092
rect 6748 20028 6749 20092
rect 6683 20027 6749 20028
rect 7419 20092 7485 20093
rect 7419 20028 7420 20092
rect 7484 20028 7485 20092
rect 7419 20027 7485 20028
rect 8155 20092 8221 20093
rect 8155 20028 8156 20092
rect 8220 20028 8221 20092
rect 8155 20027 8221 20028
rect 4865 19008 4873 19072
rect 4937 19008 4953 19072
rect 5017 19008 5033 19072
rect 5097 19008 5113 19072
rect 5177 19008 5185 19072
rect 4865 17984 5185 19008
rect 4865 17920 4873 17984
rect 4937 17920 4953 17984
rect 5017 17920 5033 17984
rect 5097 17920 5113 17984
rect 5177 17920 5185 17984
rect 4865 16896 5185 17920
rect 4865 16832 4873 16896
rect 4937 16832 4953 16896
rect 5017 16832 5033 16896
rect 5097 16832 5113 16896
rect 5177 16832 5185 16896
rect 4865 15808 5185 16832
rect 4865 15744 4873 15808
rect 4937 15744 4953 15808
rect 5017 15744 5033 15808
rect 5097 15744 5113 15808
rect 5177 15744 5185 15808
rect 4865 14720 5185 15744
rect 4865 14656 4873 14720
rect 4937 14656 4953 14720
rect 5017 14656 5033 14720
rect 5097 14656 5113 14720
rect 5177 14656 5185 14720
rect 4865 13632 5185 14656
rect 4865 13568 4873 13632
rect 4937 13568 4953 13632
rect 5017 13568 5033 13632
rect 5097 13568 5113 13632
rect 5177 13568 5185 13632
rect 4865 12544 5185 13568
rect 4865 12480 4873 12544
rect 4937 12480 4953 12544
rect 5017 12480 5033 12544
rect 5097 12480 5113 12544
rect 5177 12480 5185 12544
rect 4865 11456 5185 12480
rect 4865 11392 4873 11456
rect 4937 11392 4953 11456
rect 5017 11392 5033 11456
rect 5097 11392 5113 11456
rect 5177 11392 5185 11456
rect 4865 10368 5185 11392
rect 4865 10304 4873 10368
rect 4937 10304 4953 10368
rect 5017 10304 5033 10368
rect 5097 10304 5113 10368
rect 5177 10304 5185 10368
rect 4865 9280 5185 10304
rect 4865 9216 4873 9280
rect 4937 9216 4953 9280
rect 5017 9216 5033 9280
rect 5097 9216 5113 9280
rect 5177 9216 5185 9280
rect 4865 8192 5185 9216
rect 4865 8128 4873 8192
rect 4937 8128 4953 8192
rect 5017 8128 5033 8192
rect 5097 8128 5113 8192
rect 5177 8128 5185 8192
rect 4865 7104 5185 8128
rect 4865 7040 4873 7104
rect 4937 7040 4953 7104
rect 5017 7040 5033 7104
rect 5097 7040 5113 7104
rect 5177 7040 5185 7104
rect 4865 6016 5185 7040
rect 4865 5952 4873 6016
rect 4937 5952 4953 6016
rect 5017 5952 5033 6016
rect 5097 5952 5113 6016
rect 5177 5952 5185 6016
rect 4865 4928 5185 5952
rect 4865 4864 4873 4928
rect 4937 4864 4953 4928
rect 5017 4864 5033 4928
rect 5097 4864 5113 4928
rect 5177 4864 5185 4928
rect 4865 3840 5185 4864
rect 4865 3776 4873 3840
rect 4937 3776 4953 3840
rect 5017 3776 5033 3840
rect 5097 3776 5113 3840
rect 5177 3776 5185 3840
rect 4865 2752 5185 3776
rect 4865 2688 4873 2752
rect 4937 2688 4953 2752
rect 5017 2688 5033 2752
rect 5097 2688 5113 2752
rect 5177 2688 5185 2752
rect 4865 1664 5185 2688
rect 4865 1600 4873 1664
rect 4937 1600 4953 1664
rect 5017 1600 5033 1664
rect 5097 1600 5113 1664
rect 5177 1600 5185 1664
rect 4865 624 5185 1600
rect 8786 19616 9106 20640
rect 10366 20093 10426 21760
rect 11102 21453 11162 21760
rect 11838 21453 11898 21760
rect 11099 21452 11165 21453
rect 11099 21388 11100 21452
rect 11164 21388 11165 21452
rect 11099 21387 11165 21388
rect 11835 21452 11901 21453
rect 11835 21388 11836 21452
rect 11900 21388 11901 21452
rect 11835 21387 11901 21388
rect 12574 20365 12634 21760
rect 13310 21453 13370 21760
rect 13307 21452 13373 21453
rect 13307 21388 13308 21452
rect 13372 21388 13373 21452
rect 13307 21387 13373 21388
rect 14046 21317 14106 21760
rect 14782 21453 14842 21760
rect 15518 21453 15578 21760
rect 16254 21453 16314 21760
rect 14779 21452 14845 21453
rect 14779 21388 14780 21452
rect 14844 21388 14845 21452
rect 14779 21387 14845 21388
rect 15515 21452 15581 21453
rect 15515 21388 15516 21452
rect 15580 21388 15581 21452
rect 15515 21387 15581 21388
rect 16251 21452 16317 21453
rect 16251 21388 16252 21452
rect 16316 21388 16317 21452
rect 16251 21387 16317 21388
rect 16990 21317 17050 21760
rect 17726 21453 17786 21760
rect 18462 21453 18522 21760
rect 19198 21620 19258 21760
rect 19198 21560 19432 21620
rect 17723 21452 17789 21453
rect 17723 21388 17724 21452
rect 17788 21388 17789 21452
rect 17723 21387 17789 21388
rect 18459 21452 18525 21453
rect 18459 21388 18460 21452
rect 18524 21388 18525 21452
rect 18459 21387 18525 21388
rect 14043 21316 14109 21317
rect 14043 21252 14044 21316
rect 14108 21252 14109 21316
rect 14043 21251 14109 21252
rect 16987 21316 17053 21317
rect 16987 21252 16988 21316
rect 17052 21252 17053 21316
rect 16987 21251 17053 21252
rect 19372 21272 19432 21560
rect 19934 21453 19994 21760
rect 19931 21452 19997 21453
rect 19931 21388 19932 21452
rect 19996 21388 19997 21452
rect 19931 21387 19997 21388
rect 20300 21272 20386 21282
rect 19372 21212 20310 21272
rect 20300 21208 20310 21212
rect 20374 21208 20386 21272
rect 20300 21198 20386 21208
rect 16944 20720 17012 21178
rect 20670 20909 20730 21760
rect 21406 21453 21466 21760
rect 22142 21453 22202 21760
rect 21403 21452 21469 21453
rect 21403 21388 21404 21452
rect 21468 21388 21469 21452
rect 21403 21387 21469 21388
rect 22139 21452 22205 21453
rect 22139 21388 22140 21452
rect 22204 21388 22205 21452
rect 22139 21387 22205 21388
rect 20667 20908 20733 20909
rect 20667 20844 20668 20908
rect 20732 20844 20733 20908
rect 20667 20843 20733 20844
rect 12571 20364 12637 20365
rect 12571 20300 12572 20364
rect 12636 20300 12637 20364
rect 12571 20299 12637 20300
rect 12707 20160 13027 20720
rect 12707 20096 12715 20160
rect 12779 20096 12795 20160
rect 12859 20096 12875 20160
rect 12939 20096 12955 20160
rect 13019 20096 13027 20160
rect 10363 20092 10429 20093
rect 10363 20028 10364 20092
rect 10428 20028 10429 20092
rect 10363 20027 10429 20028
rect 8786 19552 8794 19616
rect 8858 19552 8874 19616
rect 8938 19552 8954 19616
rect 9018 19552 9034 19616
rect 9098 19552 9106 19616
rect 8786 18528 9106 19552
rect 8786 18464 8794 18528
rect 8858 18464 8874 18528
rect 8938 18464 8954 18528
rect 9018 18464 9034 18528
rect 9098 18464 9106 18528
rect 8786 17440 9106 18464
rect 8786 17376 8794 17440
rect 8858 17376 8874 17440
rect 8938 17376 8954 17440
rect 9018 17376 9034 17440
rect 9098 17376 9106 17440
rect 8786 16352 9106 17376
rect 8786 16288 8794 16352
rect 8858 16288 8874 16352
rect 8938 16288 8954 16352
rect 9018 16288 9034 16352
rect 9098 16288 9106 16352
rect 8786 15264 9106 16288
rect 8786 15200 8794 15264
rect 8858 15200 8874 15264
rect 8938 15200 8954 15264
rect 9018 15200 9034 15264
rect 9098 15200 9106 15264
rect 8786 14176 9106 15200
rect 8786 14112 8794 14176
rect 8858 14112 8874 14176
rect 8938 14112 8954 14176
rect 9018 14112 9034 14176
rect 9098 14112 9106 14176
rect 8786 13088 9106 14112
rect 8786 13024 8794 13088
rect 8858 13024 8874 13088
rect 8938 13024 8954 13088
rect 9018 13024 9034 13088
rect 9098 13024 9106 13088
rect 8786 12000 9106 13024
rect 8786 11936 8794 12000
rect 8858 11936 8874 12000
rect 8938 11936 8954 12000
rect 9018 11936 9034 12000
rect 9098 11936 9106 12000
rect 8786 10912 9106 11936
rect 8786 10848 8794 10912
rect 8858 10848 8874 10912
rect 8938 10848 8954 10912
rect 9018 10848 9034 10912
rect 9098 10848 9106 10912
rect 8786 9824 9106 10848
rect 8786 9760 8794 9824
rect 8858 9760 8874 9824
rect 8938 9760 8954 9824
rect 9018 9760 9034 9824
rect 9098 9760 9106 9824
rect 8786 8736 9106 9760
rect 8786 8672 8794 8736
rect 8858 8672 8874 8736
rect 8938 8672 8954 8736
rect 9018 8672 9034 8736
rect 9098 8672 9106 8736
rect 8786 7648 9106 8672
rect 8786 7584 8794 7648
rect 8858 7584 8874 7648
rect 8938 7584 8954 7648
rect 9018 7584 9034 7648
rect 9098 7584 9106 7648
rect 8786 6560 9106 7584
rect 8786 6496 8794 6560
rect 8858 6496 8874 6560
rect 8938 6496 8954 6560
rect 9018 6496 9034 6560
rect 9098 6496 9106 6560
rect 8786 5472 9106 6496
rect 8786 5408 8794 5472
rect 8858 5408 8874 5472
rect 8938 5408 8954 5472
rect 9018 5408 9034 5472
rect 9098 5408 9106 5472
rect 8786 4384 9106 5408
rect 8786 4320 8794 4384
rect 8858 4320 8874 4384
rect 8938 4320 8954 4384
rect 9018 4320 9034 4384
rect 9098 4320 9106 4384
rect 8786 3296 9106 4320
rect 8786 3232 8794 3296
rect 8858 3232 8874 3296
rect 8938 3232 8954 3296
rect 9018 3232 9034 3296
rect 9098 3232 9106 3296
rect 8786 2208 9106 3232
rect 8786 2144 8794 2208
rect 8858 2144 8874 2208
rect 8938 2144 8954 2208
rect 9018 2144 9034 2208
rect 9098 2144 9106 2208
rect 8786 1120 9106 2144
rect 8786 1056 8794 1120
rect 8858 1056 8874 1120
rect 8938 1056 8954 1120
rect 9018 1056 9034 1120
rect 9098 1056 9106 1120
rect 8786 1040 9106 1056
rect 12707 19072 13027 20096
rect 12707 19008 12715 19072
rect 12779 19008 12795 19072
rect 12859 19008 12875 19072
rect 12939 19008 12955 19072
rect 13019 19008 13027 19072
rect 12707 17984 13027 19008
rect 12707 17920 12715 17984
rect 12779 17920 12795 17984
rect 12859 17920 12875 17984
rect 12939 17920 12955 17984
rect 13019 17920 13027 17984
rect 12707 16896 13027 17920
rect 12707 16832 12715 16896
rect 12779 16832 12795 16896
rect 12859 16832 12875 16896
rect 12939 16832 12955 16896
rect 13019 16832 13027 16896
rect 12707 15808 13027 16832
rect 12707 15744 12715 15808
rect 12779 15744 12795 15808
rect 12859 15744 12875 15808
rect 12939 15744 12955 15808
rect 13019 15744 13027 15808
rect 12707 14720 13027 15744
rect 12707 14656 12715 14720
rect 12779 14656 12795 14720
rect 12859 14656 12875 14720
rect 12939 14656 12955 14720
rect 13019 14656 13027 14720
rect 12707 13632 13027 14656
rect 12707 13568 12715 13632
rect 12779 13568 12795 13632
rect 12859 13568 12875 13632
rect 12939 13568 12955 13632
rect 13019 13568 13027 13632
rect 12707 12544 13027 13568
rect 12707 12480 12715 12544
rect 12779 12480 12795 12544
rect 12859 12480 12875 12544
rect 12939 12480 12955 12544
rect 13019 12480 13027 12544
rect 12707 11456 13027 12480
rect 12707 11392 12715 11456
rect 12779 11392 12795 11456
rect 12859 11392 12875 11456
rect 12939 11392 12955 11456
rect 13019 11392 13027 11456
rect 12707 10368 13027 11392
rect 12707 10304 12715 10368
rect 12779 10304 12795 10368
rect 12859 10304 12875 10368
rect 12939 10304 12955 10368
rect 13019 10304 13027 10368
rect 12707 9280 13027 10304
rect 12707 9216 12715 9280
rect 12779 9216 12795 9280
rect 12859 9216 12875 9280
rect 12939 9216 12955 9280
rect 13019 9216 13027 9280
rect 12707 8192 13027 9216
rect 12707 8128 12715 8192
rect 12779 8128 12795 8192
rect 12859 8128 12875 8192
rect 12939 8128 12955 8192
rect 13019 8128 13027 8192
rect 12707 7104 13027 8128
rect 12707 7040 12715 7104
rect 12779 7040 12795 7104
rect 12859 7040 12875 7104
rect 12939 7040 12955 7104
rect 13019 7040 13027 7104
rect 12707 6016 13027 7040
rect 12707 5952 12715 6016
rect 12779 5952 12795 6016
rect 12859 5952 12875 6016
rect 12939 5952 12955 6016
rect 13019 5952 13027 6016
rect 12707 4928 13027 5952
rect 12707 4864 12715 4928
rect 12779 4864 12795 4928
rect 12859 4864 12875 4928
rect 12939 4864 12955 4928
rect 13019 4864 13027 4928
rect 12707 3840 13027 4864
rect 12707 3776 12715 3840
rect 12779 3776 12795 3840
rect 12859 3776 12875 3840
rect 12939 3776 12955 3840
rect 13019 3776 13027 3840
rect 12707 2752 13027 3776
rect 12707 2688 12715 2752
rect 12779 2688 12795 2752
rect 12859 2688 12875 2752
rect 12939 2688 12955 2752
rect 13019 2688 13027 2752
rect 12707 1664 13027 2688
rect 12707 1600 12715 1664
rect 12779 1600 12795 1664
rect 12859 1600 12875 1664
rect 12939 1600 12955 1664
rect 13019 1600 13027 1664
rect 12707 624 13027 1600
rect 16628 20704 17012 20720
rect 16628 20640 16636 20704
rect 16700 20640 16716 20704
rect 16780 20640 16796 20704
rect 16860 20640 16876 20704
rect 16940 20640 17012 20704
rect 16628 19616 17012 20640
rect 16628 19552 16636 19616
rect 16700 19552 16716 19616
rect 16780 19552 16796 19616
rect 16860 19552 16876 19616
rect 16940 19552 17012 19616
rect 16628 18528 17012 19552
rect 16628 18464 16636 18528
rect 16700 18464 16716 18528
rect 16780 18464 16796 18528
rect 16860 18464 16876 18528
rect 16940 18464 17012 18528
rect 16628 17440 17012 18464
rect 16628 17376 16636 17440
rect 16700 17376 16716 17440
rect 16780 17376 16796 17440
rect 16860 17376 16876 17440
rect 16940 17376 17012 17440
rect 16628 16352 17012 17376
rect 16628 16288 16636 16352
rect 16700 16288 16716 16352
rect 16780 16288 16796 16352
rect 16860 16288 16876 16352
rect 16940 16288 17012 16352
rect 16628 15264 17012 16288
rect 16628 15200 16636 15264
rect 16700 15200 16716 15264
rect 16780 15200 16796 15264
rect 16860 15200 16876 15264
rect 16940 15200 17012 15264
rect 16628 14176 17012 15200
rect 16628 14112 16636 14176
rect 16700 14112 16716 14176
rect 16780 14112 16796 14176
rect 16860 14112 16876 14176
rect 16940 14112 17012 14176
rect 16628 13088 17012 14112
rect 16628 13024 16636 13088
rect 16700 13024 16716 13088
rect 16780 13024 16796 13088
rect 16860 13024 16876 13088
rect 16940 13024 17012 13088
rect 16628 12000 17012 13024
rect 16628 11936 16636 12000
rect 16700 11936 16716 12000
rect 16780 11936 16796 12000
rect 16860 11936 16876 12000
rect 16940 11936 17012 12000
rect 16628 10912 17012 11936
rect 16628 10848 16636 10912
rect 16700 10848 16716 10912
rect 16780 10848 16796 10912
rect 16860 10848 16876 10912
rect 16940 10848 17012 10912
rect 16628 9824 17012 10848
rect 16628 9760 16636 9824
rect 16700 9760 16716 9824
rect 16780 9760 16796 9824
rect 16860 9760 16876 9824
rect 16940 9760 17012 9824
rect 16628 8941 17012 9760
rect 20549 20160 20869 20720
rect 22878 20501 22938 21760
rect 23614 21453 23674 21760
rect 24350 21453 24410 21760
rect 25086 21560 25146 21760
rect 25822 21453 25882 21760
rect 23611 21452 23677 21453
rect 23611 21388 23612 21452
rect 23676 21388 23677 21452
rect 23611 21387 23677 21388
rect 24347 21452 24413 21453
rect 24347 21388 24348 21452
rect 24412 21388 24413 21452
rect 24347 21387 24413 21388
rect 25819 21452 25885 21453
rect 25819 21388 25820 21452
rect 25884 21388 25885 21452
rect 25819 21387 25885 21388
rect 26558 21045 26618 21760
rect 27294 21453 27354 21760
rect 27291 21452 27357 21453
rect 27291 21388 27292 21452
rect 27356 21388 27357 21452
rect 27291 21387 27357 21388
rect 28030 21045 28090 21760
rect 28766 21453 28826 21760
rect 28763 21452 28829 21453
rect 28763 21388 28764 21452
rect 28828 21388 28829 21452
rect 28763 21387 28829 21388
rect 29502 21045 29562 21760
rect 30238 21453 30298 21760
rect 30974 21560 31034 21760
rect 31710 21560 31770 21760
rect 32446 21560 32506 21760
rect 30235 21452 30301 21453
rect 30235 21388 30236 21452
rect 30300 21388 30301 21452
rect 30235 21387 30301 21388
rect 33598 21280 33714 21294
rect 33598 21208 33614 21280
rect 33696 21230 33714 21280
rect 33696 21208 33716 21230
rect 33598 21140 33716 21208
rect 26555 21044 26621 21045
rect 26555 20980 26556 21044
rect 26620 20980 26621 21044
rect 26555 20979 26621 20980
rect 28027 21044 28093 21045
rect 28027 20980 28028 21044
rect 28092 20980 28093 21044
rect 28027 20979 28093 20980
rect 29499 21044 29565 21045
rect 29499 20980 29500 21044
rect 29564 20980 29565 21044
rect 33604 21016 33716 21140
rect 29499 20979 29565 20980
rect 24470 20704 24790 20720
rect 24470 20640 24478 20704
rect 24542 20640 24558 20704
rect 24622 20640 24638 20704
rect 24702 20640 24718 20704
rect 24782 20640 24790 20704
rect 22875 20500 22941 20501
rect 22875 20436 22876 20500
rect 22940 20436 22941 20500
rect 22875 20435 22941 20436
rect 20549 20096 20557 20160
rect 20621 20096 20637 20160
rect 20701 20096 20717 20160
rect 20781 20096 20797 20160
rect 20861 20096 20869 20160
rect 20549 19072 20869 20096
rect 20549 19008 20557 19072
rect 20621 19008 20637 19072
rect 20701 19008 20717 19072
rect 20781 19008 20797 19072
rect 20861 19008 20869 19072
rect 20549 17984 20869 19008
rect 20549 17920 20557 17984
rect 20621 17920 20637 17984
rect 20701 17920 20717 17984
rect 20781 17920 20797 17984
rect 20861 17920 20869 17984
rect 20549 16896 20869 17920
rect 20549 16832 20557 16896
rect 20621 16832 20637 16896
rect 20701 16832 20717 16896
rect 20781 16832 20797 16896
rect 20861 16832 20869 16896
rect 20549 15808 20869 16832
rect 20549 15744 20557 15808
rect 20621 15744 20637 15808
rect 20701 15744 20717 15808
rect 20781 15744 20797 15808
rect 20861 15744 20869 15808
rect 20549 14720 20869 15744
rect 20549 14656 20557 14720
rect 20621 14656 20637 14720
rect 20701 14656 20717 14720
rect 20781 14656 20797 14720
rect 20861 14656 20869 14720
rect 20549 13632 20869 14656
rect 20549 13568 20557 13632
rect 20621 13568 20637 13632
rect 20701 13568 20717 13632
rect 20781 13568 20797 13632
rect 20861 13568 20869 13632
rect 20549 12544 20869 13568
rect 20549 12480 20557 12544
rect 20621 12480 20637 12544
rect 20701 12480 20717 12544
rect 20781 12480 20797 12544
rect 20861 12480 20869 12544
rect 20549 11456 20869 12480
rect 20549 11392 20557 11456
rect 20621 11392 20637 11456
rect 20701 11392 20717 11456
rect 20781 11392 20797 11456
rect 20861 11392 20869 11456
rect 20549 10368 20869 11392
rect 20549 10304 20557 10368
rect 20621 10304 20637 10368
rect 20701 10304 20717 10368
rect 20781 10304 20797 10368
rect 20861 10304 20869 10368
rect 20549 9280 20869 10304
rect 20549 9216 20557 9280
rect 20621 9216 20637 9280
rect 20701 9216 20717 9280
rect 20781 9216 20797 9280
rect 20861 9216 20869 9280
rect 16628 8736 16948 8941
rect 16628 8672 16636 8736
rect 16700 8672 16716 8736
rect 16780 8672 16796 8736
rect 16860 8672 16876 8736
rect 16940 8672 16948 8736
rect 16628 7648 16948 8672
rect 16628 7584 16636 7648
rect 16700 7584 16716 7648
rect 16780 7584 16796 7648
rect 16860 7584 16876 7648
rect 16940 7584 16948 7648
rect 16628 6560 16948 7584
rect 16628 6496 16636 6560
rect 16700 6496 16716 6560
rect 16780 6496 16796 6560
rect 16860 6496 16876 6560
rect 16940 6496 16948 6560
rect 16628 5472 16948 6496
rect 16628 5408 16636 5472
rect 16700 5408 16716 5472
rect 16780 5408 16796 5472
rect 16860 5408 16876 5472
rect 16940 5408 16948 5472
rect 16628 4384 16948 5408
rect 16628 4320 16636 4384
rect 16700 4320 16716 4384
rect 16780 4320 16796 4384
rect 16860 4320 16876 4384
rect 16940 4320 16948 4384
rect 16628 3296 16948 4320
rect 16628 3232 16636 3296
rect 16700 3232 16716 3296
rect 16780 3232 16796 3296
rect 16860 3232 16876 3296
rect 16940 3232 16948 3296
rect 16628 2208 16948 3232
rect 16628 2144 16636 2208
rect 16700 2144 16716 2208
rect 16780 2144 16796 2208
rect 16860 2144 16876 2208
rect 16940 2144 16948 2208
rect 16628 1120 16948 2144
rect 16628 1056 16636 1120
rect 16700 1056 16716 1120
rect 16780 1056 16796 1120
rect 16860 1056 16876 1120
rect 16940 1056 16948 1120
rect 16628 1040 16948 1056
rect 20549 8192 20869 9216
rect 20549 8128 20557 8192
rect 20621 8128 20637 8192
rect 20701 8128 20717 8192
rect 20781 8128 20797 8192
rect 20861 8128 20869 8192
rect 20549 7104 20869 8128
rect 20549 7040 20557 7104
rect 20621 7040 20637 7104
rect 20701 7040 20717 7104
rect 20781 7040 20797 7104
rect 20861 7040 20869 7104
rect 20549 6016 20869 7040
rect 20549 5952 20557 6016
rect 20621 5952 20637 6016
rect 20701 5952 20717 6016
rect 20781 5952 20797 6016
rect 20861 5952 20869 6016
rect 20549 4928 20869 5952
rect 20549 4864 20557 4928
rect 20621 4864 20637 4928
rect 20701 4864 20717 4928
rect 20781 4864 20797 4928
rect 20861 4864 20869 4928
rect 20549 3840 20869 4864
rect 20549 3776 20557 3840
rect 20621 3776 20637 3840
rect 20701 3776 20717 3840
rect 20781 3776 20797 3840
rect 20861 3776 20869 3840
rect 20549 2752 20869 3776
rect 20549 2688 20557 2752
rect 20621 2688 20637 2752
rect 20701 2688 20717 2752
rect 20781 2688 20797 2752
rect 20861 2688 20869 2752
rect 20549 1664 20869 2688
rect 20549 1600 20557 1664
rect 20621 1600 20637 1664
rect 20701 1600 20717 1664
rect 20781 1600 20797 1664
rect 20861 1600 20869 1664
rect 20549 624 20869 1600
rect 24470 19616 24790 20640
rect 24470 19552 24478 19616
rect 24542 19552 24558 19616
rect 24622 19552 24638 19616
rect 24702 19552 24718 19616
rect 24782 19552 24790 19616
rect 24470 18528 24790 19552
rect 24470 18464 24478 18528
rect 24542 18464 24558 18528
rect 24622 18464 24638 18528
rect 24702 18464 24718 18528
rect 24782 18464 24790 18528
rect 24470 17440 24790 18464
rect 24470 17376 24478 17440
rect 24542 17376 24558 17440
rect 24622 17376 24638 17440
rect 24702 17376 24718 17440
rect 24782 17376 24790 17440
rect 24470 16352 24790 17376
rect 24470 16288 24478 16352
rect 24542 16288 24558 16352
rect 24622 16288 24638 16352
rect 24702 16288 24718 16352
rect 24782 16288 24790 16352
rect 24470 15264 24790 16288
rect 24470 15200 24478 15264
rect 24542 15200 24558 15264
rect 24622 15200 24638 15264
rect 24702 15200 24718 15264
rect 24782 15200 24790 15264
rect 24470 14176 24790 15200
rect 24470 14112 24478 14176
rect 24542 14112 24558 14176
rect 24622 14112 24638 14176
rect 24702 14112 24718 14176
rect 24782 14112 24790 14176
rect 24470 13088 24790 14112
rect 24470 13024 24478 13088
rect 24542 13024 24558 13088
rect 24622 13024 24638 13088
rect 24702 13024 24718 13088
rect 24782 13024 24790 13088
rect 24470 12000 24790 13024
rect 24470 11936 24478 12000
rect 24542 11936 24558 12000
rect 24622 11936 24638 12000
rect 24702 11936 24718 12000
rect 24782 11936 24790 12000
rect 24470 10912 24790 11936
rect 24470 10848 24478 10912
rect 24542 10848 24558 10912
rect 24622 10848 24638 10912
rect 24702 10848 24718 10912
rect 24782 10848 24790 10912
rect 24470 9824 24790 10848
rect 24470 9760 24478 9824
rect 24542 9760 24558 9824
rect 24622 9760 24638 9824
rect 24702 9760 24718 9824
rect 24782 9760 24790 9824
rect 24470 8736 24790 9760
rect 24470 8672 24478 8736
rect 24542 8672 24558 8736
rect 24622 8672 24638 8736
rect 24702 8672 24718 8736
rect 24782 8672 24790 8736
rect 24470 7648 24790 8672
rect 24470 7584 24478 7648
rect 24542 7584 24558 7648
rect 24622 7584 24638 7648
rect 24702 7584 24718 7648
rect 24782 7584 24790 7648
rect 24470 6560 24790 7584
rect 24470 6496 24478 6560
rect 24542 6496 24558 6560
rect 24622 6496 24638 6560
rect 24702 6496 24718 6560
rect 24782 6496 24790 6560
rect 24470 5472 24790 6496
rect 24470 5408 24478 5472
rect 24542 5408 24558 5472
rect 24622 5408 24638 5472
rect 24702 5408 24718 5472
rect 24782 5408 24790 5472
rect 24470 4384 24790 5408
rect 24470 4320 24478 4384
rect 24542 4320 24558 4384
rect 24622 4320 24638 4384
rect 24702 4320 24718 4384
rect 24782 4320 24790 4384
rect 24470 3296 24790 4320
rect 24470 3232 24478 3296
rect 24542 3232 24558 3296
rect 24622 3232 24638 3296
rect 24702 3232 24718 3296
rect 24782 3232 24790 3296
rect 24470 2208 24790 3232
rect 24470 2144 24478 2208
rect 24542 2144 24558 2208
rect 24622 2144 24638 2208
rect 24702 2144 24718 2208
rect 24782 2144 24790 2208
rect 24470 1120 24790 2144
rect 24470 1056 24478 1120
rect 24542 1056 24558 1120
rect 24622 1056 24638 1120
rect 24702 1056 24718 1120
rect 24782 1056 24790 1120
rect 24470 1040 24790 1056
rect 28391 20160 28711 20720
rect 28391 20096 28399 20160
rect 28463 20096 28479 20160
rect 28543 20096 28559 20160
rect 28623 20096 28639 20160
rect 28703 20096 28711 20160
rect 28391 19072 28711 20096
rect 28391 19008 28399 19072
rect 28463 19008 28479 19072
rect 28543 19008 28559 19072
rect 28623 19008 28639 19072
rect 28703 19008 28711 19072
rect 28391 17984 28711 19008
rect 28391 17920 28399 17984
rect 28463 17920 28479 17984
rect 28543 17920 28559 17984
rect 28623 17920 28639 17984
rect 28703 17920 28711 17984
rect 28391 16896 28711 17920
rect 28391 16832 28399 16896
rect 28463 16832 28479 16896
rect 28543 16832 28559 16896
rect 28623 16832 28639 16896
rect 28703 16832 28711 16896
rect 28391 15808 28711 16832
rect 28391 15744 28399 15808
rect 28463 15744 28479 15808
rect 28543 15744 28559 15808
rect 28623 15744 28639 15808
rect 28703 15744 28711 15808
rect 28391 14720 28711 15744
rect 28391 14656 28399 14720
rect 28463 14656 28479 14720
rect 28543 14656 28559 14720
rect 28623 14656 28639 14720
rect 28703 14656 28711 14720
rect 28391 13632 28711 14656
rect 28391 13568 28399 13632
rect 28463 13568 28479 13632
rect 28543 13568 28559 13632
rect 28623 13568 28639 13632
rect 28703 13568 28711 13632
rect 28391 12544 28711 13568
rect 28391 12480 28399 12544
rect 28463 12480 28479 12544
rect 28543 12480 28559 12544
rect 28623 12480 28639 12544
rect 28703 12480 28711 12544
rect 28391 11456 28711 12480
rect 28391 11392 28399 11456
rect 28463 11392 28479 11456
rect 28543 11392 28559 11456
rect 28623 11392 28639 11456
rect 28703 11392 28711 11456
rect 28391 10368 28711 11392
rect 28391 10304 28399 10368
rect 28463 10304 28479 10368
rect 28543 10304 28559 10368
rect 28623 10304 28639 10368
rect 28703 10304 28711 10368
rect 28391 9280 28711 10304
rect 28391 9216 28399 9280
rect 28463 9216 28479 9280
rect 28543 9216 28559 9280
rect 28623 9216 28639 9280
rect 28703 9216 28711 9280
rect 28391 8192 28711 9216
rect 28391 8128 28399 8192
rect 28463 8128 28479 8192
rect 28543 8128 28559 8192
rect 28623 8128 28639 8192
rect 28703 8128 28711 8192
rect 28391 7104 28711 8128
rect 28391 7040 28399 7104
rect 28463 7040 28479 7104
rect 28543 7040 28559 7104
rect 28623 7040 28639 7104
rect 28703 7040 28711 7104
rect 28391 6016 28711 7040
rect 28391 5952 28399 6016
rect 28463 5952 28479 6016
rect 28543 5952 28559 6016
rect 28623 5952 28639 6016
rect 28703 5952 28711 6016
rect 28391 4928 28711 5952
rect 28391 4864 28399 4928
rect 28463 4864 28479 4928
rect 28543 4864 28559 4928
rect 28623 4864 28639 4928
rect 28703 4864 28711 4928
rect 28391 3840 28711 4864
rect 28391 3776 28399 3840
rect 28463 3776 28479 3840
rect 28543 3776 28559 3840
rect 28623 3776 28639 3840
rect 28703 3776 28711 3840
rect 28391 2752 28711 3776
rect 28391 2688 28399 2752
rect 28463 2688 28479 2752
rect 28543 2688 28559 2752
rect 28623 2688 28639 2752
rect 28703 2688 28711 2752
rect 28391 1664 28711 2688
rect 28391 1600 28399 1664
rect 28463 1600 28479 1664
rect 28543 1600 28559 1664
rect 28623 1600 28639 1664
rect 28703 1600 28711 1664
rect 28391 624 28711 1600
rect 32312 20704 32632 20720
rect 32312 20640 32320 20704
rect 32384 20640 32400 20704
rect 32464 20640 32480 20704
rect 32544 20640 32560 20704
rect 32624 20640 32632 20704
rect 32312 19616 32632 20640
rect 32312 19552 32320 19616
rect 32384 19552 32400 19616
rect 32464 19552 32480 19616
rect 32544 19552 32560 19616
rect 32624 19552 32632 19616
rect 32312 18528 32632 19552
rect 32312 18464 32320 18528
rect 32384 18464 32400 18528
rect 32464 18464 32480 18528
rect 32544 18464 32560 18528
rect 32624 18464 32632 18528
rect 32312 17440 32632 18464
rect 32312 17376 32320 17440
rect 32384 17376 32400 17440
rect 32464 17376 32480 17440
rect 32544 17376 32560 17440
rect 32624 17376 32632 17440
rect 32312 16352 32632 17376
rect 32312 16288 32320 16352
rect 32384 16288 32400 16352
rect 32464 16288 32480 16352
rect 32544 16288 32560 16352
rect 32624 16288 32632 16352
rect 32312 15264 32632 16288
rect 32312 15200 32320 15264
rect 32384 15200 32400 15264
rect 32464 15200 32480 15264
rect 32544 15200 32560 15264
rect 32624 15200 32632 15264
rect 32312 14176 32632 15200
rect 32312 14112 32320 14176
rect 32384 14112 32400 14176
rect 32464 14112 32480 14176
rect 32544 14112 32560 14176
rect 32624 14112 32632 14176
rect 32312 13088 32632 14112
rect 32312 13024 32320 13088
rect 32384 13024 32400 13088
rect 32464 13024 32480 13088
rect 32544 13024 32560 13088
rect 32624 13024 32632 13088
rect 32312 12000 32632 13024
rect 32312 11936 32320 12000
rect 32384 11936 32400 12000
rect 32464 11936 32480 12000
rect 32544 11936 32560 12000
rect 32624 11936 32632 12000
rect 32312 10912 32632 11936
rect 32312 10848 32320 10912
rect 32384 10848 32400 10912
rect 32464 10848 32480 10912
rect 32544 10848 32560 10912
rect 32624 10848 32632 10912
rect 32312 9824 32632 10848
rect 32312 9760 32320 9824
rect 32384 9760 32400 9824
rect 32464 9760 32480 9824
rect 32544 9760 32560 9824
rect 32624 9760 32632 9824
rect 32312 8736 32632 9760
rect 32312 8672 32320 8736
rect 32384 8672 32400 8736
rect 32464 8672 32480 8736
rect 32544 8672 32560 8736
rect 32624 8672 32632 8736
rect 32312 7648 32632 8672
rect 32312 7584 32320 7648
rect 32384 7584 32400 7648
rect 32464 7584 32480 7648
rect 32544 7584 32560 7648
rect 32624 7584 32632 7648
rect 32312 6560 32632 7584
rect 32312 6496 32320 6560
rect 32384 6496 32400 6560
rect 32464 6496 32480 6560
rect 32544 6496 32560 6560
rect 32624 6496 32632 6560
rect 32312 5472 32632 6496
rect 32312 5408 32320 5472
rect 32384 5408 32400 5472
rect 32464 5408 32480 5472
rect 32544 5408 32560 5472
rect 32624 5408 32632 5472
rect 32312 4384 32632 5408
rect 32312 4320 32320 4384
rect 32384 4320 32400 4384
rect 32464 4320 32480 4384
rect 32544 4320 32560 4384
rect 32624 4320 32632 4384
rect 32312 3296 32632 4320
rect 32312 3232 32320 3296
rect 32384 3232 32400 3296
rect 32464 3232 32480 3296
rect 32544 3232 32560 3296
rect 32624 3232 32632 3296
rect 32312 2208 32632 3232
rect 32312 2144 32320 2208
rect 32384 2144 32400 2208
rect 32464 2144 32480 2208
rect 32544 2144 32560 2208
rect 32624 2144 32632 2208
rect 32312 1120 32632 2144
rect 32312 1056 32320 1120
rect 32384 1056 32400 1120
rect 32464 1056 32480 1120
rect 32544 1056 32560 1120
rect 32624 1056 32632 1120
rect -54 266 2602 320
rect 4865 304 28716 624
rect -54 -330 2890 266
rect -52 -408 2890 -330
rect 2132 -605 2890 -408
rect 2132 -634 13797 -605
rect 2132 -882 2172 -634
rect 13766 -882 13797 -634
rect 2132 -907 13797 -882
rect 15882 -2320 16202 304
rect 32312 -140 32632 1056
rect 2120 -2342 16202 -2320
rect 1058 -2470 1568 -2446
rect 1058 -2636 1262 -2470
rect 1526 -2636 1568 -2470
rect 1058 -3032 1568 -2636
rect 2120 -2598 2134 -2342
rect 13776 -2598 16202 -2342
rect 2120 -2640 16202 -2598
rect 18530 -460 32632 -140
rect 1158 -4278 1274 -3032
rect 18530 -3178 18850 -460
rect 20268 -1705 20384 -1702
rect 33605 -1705 33715 21016
rect 20268 -1815 33715 -1705
rect 18252 -3302 18956 -3178
rect 18252 -3734 18388 -3302
rect 18836 -3734 18956 -3302
rect 18252 -3810 18956 -3734
rect 20268 -4278 20384 -1815
rect 1158 -4394 20384 -4278
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1685868990
transform 1 0 2484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1685868990
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1685868990
transform 1 0 4876 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1685868990
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1685868990
transform 1 0 7452 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1685868990
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1685868990
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1685868990
transform 1 0 10028 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1685868990
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1685868990
transform 1 0 11500 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1685868990
transform 1 0 12604 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1685868990
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1685868990
transform 1 0 14076 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1685868990
transform 1 0 15180 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1685868990
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1685868990
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1685868990
transform 1 0 17756 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1685868990
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1685868990
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1685868990
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1685868990
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1685868990
transform 1 0 21804 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1685868990
transform 1 0 22908 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1685868990
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1685868990
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1685868990
transform 1 0 25484 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1685868990
transform 1 0 26588 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1685868990
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1685868990
transform 1 0 28060 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1685868990
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1685868990
transform 1 0 29532 0 1 1088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1685868990
transform 1 0 30636 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1685868990
transform 1 0 31740 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_337
timestamp 1685868990
transform 1 0 32108 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1685868990
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1685868990
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1685868990
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1685868990
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1685868990
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1685868990
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1685868990
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1685868990
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1685868990
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1685868990
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1685868990
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1685868990
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1685868990
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1685868990
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1685868990
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1685868990
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1685868990
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1685868990
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1685868990
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1685868990
transform 1 0 19964 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1685868990
transform 1 0 21068 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1685868990
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1685868990
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1685868990
transform 1 0 22908 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1685868990
transform 1 0 24012 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1685868990
transform 1 0 25116 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1685868990
transform 1 0 26220 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1685868990
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1685868990
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1685868990
transform 1 0 28060 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1685868990
transform 1 0 29164 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1685868990
transform 1 0 30268 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1685868990
transform 1 0 31372 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1685868990
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_337
timestamp 1685868990
transform 1 0 32108 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1685868990
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1685868990
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1685868990
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1685868990
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1685868990
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1685868990
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1685868990
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1685868990
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1685868990
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1685868990
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1685868990
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1685868990
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1685868990
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1685868990
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1685868990
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1685868990
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1685868990
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1685868990
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1685868990
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1685868990
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1685868990
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1685868990
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1685868990
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1685868990
transform 1 0 21436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1685868990
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1685868990
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1685868990
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1685868990
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1685868990
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1685868990
transform 1 0 26588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1685868990
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1685868990
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1685868990
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1685868990
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1685868990
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_333
timestamp 1685868990
transform 1 0 31740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_337
timestamp 1685868990
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1685868990
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1685868990
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1685868990
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1685868990
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1685868990
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1685868990
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1685868990
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1685868990
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1685868990
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1685868990
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1685868990
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1685868990
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1685868990
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1685868990
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1685868990
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1685868990
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1685868990
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1685868990
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1685868990
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1685868990
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1685868990
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1685868990
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1685868990
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1685868990
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1685868990
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1685868990
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1685868990
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1685868990
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1685868990
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1685868990
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1685868990
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1685868990
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1685868990
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1685868990
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1685868990
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1685868990
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp 1685868990
transform 1 0 32108 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1685868990
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1685868990
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1685868990
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1685868990
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1685868990
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1685868990
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1685868990
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1685868990
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1685868990
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1685868990
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1685868990
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1685868990
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1685868990
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1685868990
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1685868990
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1685868990
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1685868990
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1685868990
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1685868990
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1685868990
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1685868990
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1685868990
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1685868990
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1685868990
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1685868990
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1685868990
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1685868990
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1685868990
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1685868990
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1685868990
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1685868990
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1685868990
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1685868990
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1685868990
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1685868990
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_333
timestamp 1685868990
transform 1 0 31740 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_337
timestamp 1685868990
transform 1 0 32108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1685868990
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1685868990
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1685868990
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1685868990
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1685868990
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1685868990
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1685868990
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1685868990
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1685868990
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1685868990
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1685868990
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1685868990
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1685868990
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1685868990
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1685868990
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1685868990
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1685868990
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1685868990
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1685868990
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1685868990
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1685868990
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1685868990
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1685868990
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1685868990
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1685868990
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1685868990
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1685868990
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1685868990
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1685868990
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1685868990
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1685868990
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1685868990
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1685868990
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1685868990
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1685868990
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1685868990
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_337
timestamp 1685868990
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1685868990
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1685868990
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1685868990
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1685868990
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1685868990
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1685868990
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1685868990
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1685868990
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1685868990
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1685868990
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1685868990
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1685868990
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1685868990
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1685868990
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1685868990
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1685868990
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1685868990
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1685868990
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1685868990
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1685868990
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1685868990
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1685868990
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1685868990
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1685868990
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1685868990
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1685868990
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1685868990
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1685868990
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1685868990
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1685868990
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1685868990
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1685868990
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1685868990
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1685868990
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1685868990
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_333
timestamp 1685868990
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_337
timestamp 1685868990
transform 1 0 32108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1685868990
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1685868990
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1685868990
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1685868990
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1685868990
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1685868990
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1685868990
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1685868990
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1685868990
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1685868990
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1685868990
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1685868990
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1685868990
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1685868990
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1685868990
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1685868990
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1685868990
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1685868990
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1685868990
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1685868990
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1685868990
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1685868990
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1685868990
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1685868990
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1685868990
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1685868990
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1685868990
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1685868990
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1685868990
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1685868990
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1685868990
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1685868990
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1685868990
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1685868990
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1685868990
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1685868990
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_337
timestamp 1685868990
transform 1 0 32108 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1685868990
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1685868990
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1685868990
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1685868990
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1685868990
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1685868990
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1685868990
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1685868990
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1685868990
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1685868990
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1685868990
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1685868990
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1685868990
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1685868990
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1685868990
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1685868990
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1685868990
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1685868990
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1685868990
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1685868990
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1685868990
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1685868990
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1685868990
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1685868990
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1685868990
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1685868990
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1685868990
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1685868990
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1685868990
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1685868990
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1685868990
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1685868990
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1685868990
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1685868990
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1685868990
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_333
timestamp 1685868990
transform 1 0 31740 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_337
timestamp 1685868990
transform 1 0 32108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1685868990
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1685868990
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1685868990
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1685868990
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1685868990
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1685868990
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1685868990
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1685868990
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1685868990
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1685868990
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1685868990
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1685868990
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1685868990
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1685868990
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1685868990
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1685868990
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1685868990
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1685868990
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1685868990
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1685868990
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1685868990
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1685868990
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1685868990
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1685868990
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1685868990
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1685868990
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1685868990
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1685868990
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1685868990
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1685868990
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1685868990
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1685868990
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1685868990
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1685868990
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1685868990
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1685868990
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_337
timestamp 1685868990
transform 1 0 32108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1685868990
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1685868990
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1685868990
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1685868990
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1685868990
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1685868990
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1685868990
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1685868990
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1685868990
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1685868990
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1685868990
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1685868990
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1685868990
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1685868990
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1685868990
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1685868990
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1685868990
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1685868990
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1685868990
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1685868990
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1685868990
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1685868990
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1685868990
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1685868990
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1685868990
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1685868990
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1685868990
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1685868990
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1685868990
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1685868990
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1685868990
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1685868990
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1685868990
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1685868990
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1685868990
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_333
timestamp 1685868990
transform 1 0 31740 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_337
timestamp 1685868990
transform 1 0 32108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1685868990
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1685868990
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1685868990
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1685868990
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1685868990
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1685868990
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1685868990
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1685868990
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1685868990
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1685868990
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1685868990
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1685868990
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1685868990
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1685868990
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1685868990
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1685868990
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1685868990
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1685868990
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1685868990
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1685868990
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1685868990
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1685868990
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1685868990
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1685868990
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1685868990
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1685868990
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1685868990
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1685868990
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1685868990
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1685868990
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1685868990
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1685868990
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1685868990
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1685868990
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1685868990
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1685868990
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_337
timestamp 1685868990
transform 1 0 32108 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1685868990
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1685868990
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1685868990
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1685868990
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1685868990
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1685868990
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1685868990
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1685868990
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1685868990
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1685868990
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1685868990
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1685868990
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1685868990
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1685868990
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1685868990
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1685868990
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1685868990
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1685868990
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1685868990
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1685868990
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1685868990
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1685868990
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1685868990
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1685868990
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1685868990
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1685868990
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1685868990
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1685868990
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1685868990
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1685868990
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1685868990
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1685868990
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1685868990
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1685868990
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1685868990
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1685868990
transform 1 0 31740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_337
timestamp 1685868990
transform 1 0 32108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1685868990
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1685868990
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1685868990
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1685868990
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1685868990
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1685868990
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1685868990
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1685868990
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1685868990
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1685868990
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1685868990
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1685868990
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1685868990
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1685868990
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1685868990
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1685868990
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1685868990
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1685868990
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1685868990
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1685868990
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1685868990
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1685868990
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1685868990
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1685868990
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1685868990
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1685868990
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1685868990
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1685868990
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1685868990
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1685868990
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1685868990
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1685868990
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1685868990
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1685868990
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1685868990
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1685868990
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_337
timestamp 1685868990
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1685868990
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1685868990
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1685868990
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1685868990
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1685868990
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1685868990
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1685868990
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1685868990
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1685868990
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1685868990
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1685868990
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1685868990
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1685868990
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1685868990
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1685868990
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1685868990
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1685868990
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1685868990
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1685868990
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1685868990
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1685868990
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1685868990
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1685868990
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1685868990
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1685868990
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1685868990
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1685868990
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1685868990
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1685868990
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1685868990
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1685868990
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1685868990
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1685868990
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1685868990
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1685868990
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_333
timestamp 1685868990
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_337
timestamp 1685868990
transform 1 0 32108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1685868990
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1685868990
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1685868990
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1685868990
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1685868990
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1685868990
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1685868990
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1685868990
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1685868990
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1685868990
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1685868990
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1685868990
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1685868990
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1685868990
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1685868990
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1685868990
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1685868990
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1685868990
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1685868990
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1685868990
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1685868990
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1685868990
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1685868990
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1685868990
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1685868990
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1685868990
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1685868990
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1685868990
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1685868990
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1685868990
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1685868990
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1685868990
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1685868990
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1685868990
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1685868990
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1685868990
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_337
timestamp 1685868990
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1685868990
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1685868990
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1685868990
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1685868990
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1685868990
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1685868990
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1685868990
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1685868990
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1685868990
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1685868990
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1685868990
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1685868990
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1685868990
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1685868990
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1685868990
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1685868990
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1685868990
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1685868990
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1685868990
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1685868990
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1685868990
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1685868990
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1685868990
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1685868990
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1685868990
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1685868990
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1685868990
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1685868990
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1685868990
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1685868990
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1685868990
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1685868990
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1685868990
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1685868990
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1685868990
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_333
timestamp 1685868990
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_337
timestamp 1685868990
transform 1 0 32108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1685868990
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1685868990
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1685868990
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1685868990
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1685868990
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1685868990
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1685868990
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1685868990
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1685868990
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1685868990
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1685868990
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1685868990
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1685868990
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1685868990
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1685868990
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1685868990
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1685868990
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1685868990
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1685868990
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1685868990
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1685868990
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1685868990
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1685868990
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1685868990
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1685868990
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1685868990
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1685868990
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1685868990
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1685868990
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1685868990
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1685868990
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1685868990
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1685868990
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1685868990
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1685868990
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1685868990
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_337
timestamp 1685868990
transform 1 0 32108 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1685868990
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1685868990
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1685868990
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1685868990
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1685868990
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1685868990
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1685868990
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1685868990
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1685868990
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1685868990
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1685868990
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1685868990
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1685868990
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1685868990
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1685868990
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1685868990
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1685868990
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1685868990
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1685868990
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1685868990
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1685868990
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1685868990
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1685868990
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1685868990
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1685868990
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1685868990
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1685868990
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1685868990
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1685868990
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1685868990
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1685868990
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1685868990
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1685868990
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1685868990
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1685868990
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_333
timestamp 1685868990
transform 1 0 31740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_337
timestamp 1685868990
transform 1 0 32108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1685868990
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1685868990
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1685868990
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1685868990
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1685868990
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1685868990
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1685868990
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1685868990
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1685868990
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1685868990
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1685868990
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1685868990
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1685868990
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1685868990
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1685868990
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1685868990
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1685868990
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1685868990
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1685868990
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1685868990
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1685868990
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1685868990
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1685868990
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1685868990
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1685868990
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1685868990
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1685868990
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1685868990
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1685868990
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1685868990
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1685868990
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1685868990
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1685868990
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1685868990
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1685868990
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1685868990
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_337
timestamp 1685868990
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1685868990
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1685868990
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1685868990
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1685868990
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1685868990
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1685868990
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1685868990
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1685868990
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1685868990
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1685868990
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1685868990
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1685868990
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1685868990
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1685868990
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1685868990
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1685868990
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1685868990
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1685868990
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1685868990
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1685868990
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1685868990
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1685868990
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1685868990
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1685868990
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_228
timestamp 1685868990
transform 1 0 22080 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1685868990
transform 1 0 23184 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1685868990
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1685868990
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1685868990
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1685868990
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1685868990
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1685868990
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1685868990
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1685868990
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_333
timestamp 1685868990
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_337
timestamp 1685868990
transform 1 0 32108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1685868990
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1685868990
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1685868990
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1685868990
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1685868990
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1685868990
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1685868990
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1685868990
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1685868990
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1685868990
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1685868990
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1685868990
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1685868990
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1685868990
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1685868990
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1685868990
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1685868990
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1685868990
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1685868990
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1685868990
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1685868990
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1685868990
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1685868990
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1685868990
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1685868990
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_237 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 23644 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_254
timestamp 1685868990
transform 1 0 24472 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_266
timestamp 1685868990
transform 1 0 25576 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1685868990
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1685868990
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1685868990
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1685868990
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1685868990
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1685868990
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1685868990
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_337
timestamp 1685868990
transform 1 0 32108 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1685868990
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1685868990
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1685868990
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1685868990
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1685868990
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1685868990
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1685868990
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1685868990
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1685868990
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1685868990
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1685868990
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1685868990
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1685868990
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1685868990
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1685868990
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1685868990
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1685868990
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1685868990
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1685868990
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1685868990
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1685868990
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1685868990
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1685868990
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1685868990
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1685868990
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1685868990
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1685868990
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1685868990
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1685868990
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1685868990
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1685868990
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1685868990
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1685868990
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1685868990
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1685868990
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_333
timestamp 1685868990
transform 1 0 31740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_337
timestamp 1685868990
transform 1 0 32108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1685868990
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1685868990
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1685868990
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1685868990
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1685868990
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1685868990
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1685868990
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1685868990
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1685868990
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1685868990
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1685868990
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1685868990
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1685868990
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1685868990
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1685868990
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1685868990
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1685868990
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1685868990
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1685868990
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1685868990
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1685868990
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1685868990
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1685868990
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1685868990
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1685868990
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1685868990
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_249
timestamp 1685868990
transform 1 0 24012 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_255
timestamp 1685868990
transform 1 0 24564 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1685868990
transform 1 0 25116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_270
timestamp 1685868990
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1685868990
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1685868990
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1685868990
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1685868990
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1685868990
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1685868990
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1685868990
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_337
timestamp 1685868990
transform 1 0 32108 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1685868990
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1685868990
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1685868990
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1685868990
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1685868990
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1685868990
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1685868990
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1685868990
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1685868990
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1685868990
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1685868990
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1685868990
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1685868990
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1685868990
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1685868990
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1685868990
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1685868990
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1685868990
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1685868990
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1685868990
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1685868990
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_197
timestamp 1685868990
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1685868990
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_212
timestamp 1685868990
transform 1 0 20608 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_224
timestamp 1685868990
transform 1 0 21712 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_236
timestamp 1685868990
transform 1 0 22816 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1685868990
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1685868990
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1685868990
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1685868990
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1685868990
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1685868990
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1685868990
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1685868990
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1685868990
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_333
timestamp 1685868990
transform 1 0 31740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_337
timestamp 1685868990
transform 1 0 32108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1685868990
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1685868990
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1685868990
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1685868990
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1685868990
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1685868990
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1685868990
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1685868990
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1685868990
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1685868990
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1685868990
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1685868990
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1685868990
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1685868990
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1685868990
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1685868990
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1685868990
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1685868990
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1685868990
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1685868990
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1685868990
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1685868990
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1685868990
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1685868990
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1685868990
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1685868990
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_249
timestamp 1685868990
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_255
timestamp 1685868990
transform 1 0 24564 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_266
timestamp 1685868990
transform 1 0 25576 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1685868990
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1685868990
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1685868990
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1685868990
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1685868990
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1685868990
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1685868990
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_337
timestamp 1685868990
transform 1 0 32108 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1685868990
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1685868990
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1685868990
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1685868990
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1685868990
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1685868990
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1685868990
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1685868990
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1685868990
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1685868990
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1685868990
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1685868990
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1685868990
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1685868990
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1685868990
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1685868990
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1685868990
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1685868990
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1685868990
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1685868990
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1685868990
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1685868990
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1685868990
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1685868990
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1685868990
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1685868990
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1685868990
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1685868990
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1685868990
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1685868990
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1685868990
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1685868990
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1685868990
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1685868990
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1685868990
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_333
timestamp 1685868990
transform 1 0 31740 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_337
timestamp 1685868990
transform 1 0 32108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1685868990
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1685868990
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1685868990
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1685868990
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1685868990
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1685868990
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1685868990
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1685868990
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1685868990
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1685868990
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1685868990
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1685868990
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1685868990
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1685868990
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1685868990
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1685868990
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1685868990
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1685868990
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1685868990
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_187
timestamp 1685868990
transform 1 0 18308 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_199
timestamp 1685868990
transform 1 0 19412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_211
timestamp 1685868990
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1685868990
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1685868990
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1685868990
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1685868990
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1685868990
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1685868990
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1685868990
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1685868990
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1685868990
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1685868990
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1685868990
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1685868990
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1685868990
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_337
timestamp 1685868990
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1685868990
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1685868990
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1685868990
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1685868990
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1685868990
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1685868990
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1685868990
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1685868990
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1685868990
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1685868990
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1685868990
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1685868990
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1685868990
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1685868990
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1685868990
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1685868990
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1685868990
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1685868990
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1685868990
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1685868990
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1685868990
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1685868990
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1685868990
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1685868990
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_233
timestamp 1685868990
transform 1 0 22540 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_239
timestamp 1685868990
transform 1 0 23092 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1685868990
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1685868990
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 1685868990
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_258
timestamp 1685868990
transform 1 0 24840 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_270
timestamp 1685868990
transform 1 0 25944 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_282
timestamp 1685868990
transform 1 0 27048 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_294
timestamp 1685868990
transform 1 0 28152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1685868990
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1685868990
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1685868990
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_333
timestamp 1685868990
transform 1 0 31740 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_337
timestamp 1685868990
transform 1 0 32108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1685868990
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1685868990
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1685868990
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1685868990
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1685868990
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1685868990
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1685868990
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1685868990
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1685868990
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1685868990
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1685868990
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1685868990
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1685868990
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1685868990
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1685868990
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1685868990
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1685868990
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1685868990
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1685868990
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1685868990
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1685868990
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1685868990
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1685868990
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1685868990
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1685868990
transform 1 0 21804 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_248
timestamp 1685868990
transform 1 0 23920 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_260
timestamp 1685868990
transform 1 0 25024 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1685868990
transform 1 0 26128 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1685868990
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1685868990
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1685868990
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1685868990
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1685868990
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1685868990
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_337
timestamp 1685868990
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1685868990
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1685868990
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1685868990
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1685868990
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1685868990
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1685868990
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1685868990
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1685868990
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1685868990
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1685868990
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1685868990
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1685868990
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1685868990
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1685868990
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1685868990
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1685868990
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1685868990
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1685868990
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1685868990
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1685868990
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1685868990
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1685868990
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1685868990
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1685868990
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_233
timestamp 1685868990
transform 1 0 22540 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_241
timestamp 1685868990
transform 1 0 23276 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1685868990
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1685868990
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1685868990
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1685868990
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1685868990
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1685868990
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1685868990
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1685868990
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1685868990
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1685868990
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_333
timestamp 1685868990
transform 1 0 31740 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_337
timestamp 1685868990
transform 1 0 32108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1685868990
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1685868990
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1685868990
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1685868990
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1685868990
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1685868990
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1685868990
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1685868990
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1685868990
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1685868990
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1685868990
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1685868990
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1685868990
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1685868990
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1685868990
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1685868990
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1685868990
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1685868990
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1685868990
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1685868990
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1685868990
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1685868990
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1685868990
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1685868990
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1685868990
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_237
timestamp 1685868990
transform 1 0 22908 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_246
timestamp 1685868990
transform 1 0 23736 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_258
timestamp 1685868990
transform 1 0 24840 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_270
timestamp 1685868990
transform 1 0 25944 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1685868990
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1685868990
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1685868990
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1685868990
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1685868990
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1685868990
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1685868990
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_337
timestamp 1685868990
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1685868990
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1685868990
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1685868990
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1685868990
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1685868990
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1685868990
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1685868990
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1685868990
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1685868990
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1685868990
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1685868990
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1685868990
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1685868990
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1685868990
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1685868990
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1685868990
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_175
timestamp 1685868990
transform 1 0 17204 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_179
timestamp 1685868990
transform 1 0 17572 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1685868990
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1685868990
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1685868990
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1685868990
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_221
timestamp 1685868990
transform 1 0 21436 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_227
timestamp 1685868990
transform 1 0 21988 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_231
timestamp 1685868990
transform 1 0 22356 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_238
timestamp 1685868990
transform 1 0 23000 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1685868990
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_253
timestamp 1685868990
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_262
timestamp 1685868990
transform 1 0 25208 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_274
timestamp 1685868990
transform 1 0 26312 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_286
timestamp 1685868990
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1685868990
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1685868990
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1685868990
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1685868990
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1685868990
transform 1 0 31740 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_337
timestamp 1685868990
transform 1 0 32108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1685868990
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1685868990
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1685868990
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1685868990
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1685868990
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1685868990
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1685868990
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1685868990
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_81
timestamp 1685868990
transform 1 0 8556 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_88
timestamp 1685868990
transform 1 0 9200 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_100
timestamp 1685868990
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1685868990
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_120
timestamp 1685868990
transform 1 0 12144 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_132
timestamp 1685868990
transform 1 0 13248 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_144
timestamp 1685868990
transform 1 0 14352 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_156
timestamp 1685868990
transform 1 0 15456 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1685868990
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1685868990
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_201
timestamp 1685868990
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_207
timestamp 1685868990
transform 1 0 20148 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1685868990
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1685868990
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_230
timestamp 1685868990
transform 1 0 22264 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_241
timestamp 1685868990
transform 1 0 23276 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_249
timestamp 1685868990
transform 1 0 24012 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_257
timestamp 1685868990
transform 1 0 24748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1685868990
transform 1 0 25852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1685868990
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1685868990
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1685868990
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1685868990
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1685868990
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1685868990
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1685868990
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_337
timestamp 1685868990
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1685868990
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1685868990
transform 1 0 1840 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1685868990
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1685868990
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1685868990
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_53
timestamp 1685868990
transform 1 0 5980 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1685868990
transform 1 0 6992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_68
timestamp 1685868990
transform 1 0 7360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_72
timestamp 1685868990
transform 1 0 7728 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_76
timestamp 1685868990
transform 1 0 8096 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1685868990
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1685868990
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1685868990
transform 1 0 9568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1685868990
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_106
timestamp 1685868990
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1685868990
transform 1 0 11684 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_123
timestamp 1685868990
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1685868990
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1685868990
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1685868990
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1685868990
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1685868990
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_177
timestamp 1685868990
transform 1 0 17388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_186
timestamp 1685868990
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1685868990
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1685868990
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_204
timestamp 1685868990
transform 1 0 19872 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_212
timestamp 1685868990
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_217
timestamp 1685868990
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_226
timestamp 1685868990
transform 1 0 21896 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1685868990
transform 1 0 22724 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1685868990
transform 1 0 23552 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1685868990
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1685868990
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1685868990
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1685868990
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1685868990
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1685868990
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1685868990
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1685868990
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1685868990
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_337
timestamp 1685868990
transform 1 0 32108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1685868990
transform 1 0 1380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_12
timestamp 1685868990
transform 1 0 2208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_19
timestamp 1685868990
transform 1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_26
timestamp 1685868990
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_29
timestamp 1685868990
transform 1 0 3772 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_40
timestamp 1685868990
transform 1 0 4784 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_47
timestamp 1685868990
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1685868990
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1685868990
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_81
timestamp 1685868990
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_85
timestamp 1685868990
transform 1 0 8924 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_91
timestamp 1685868990
transform 1 0 9476 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_107
timestamp 1685868990
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1685868990
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_113
timestamp 1685868990
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_138
timestamp 1685868990
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_141
timestamp 1685868990
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_153
timestamp 1685868990
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1685868990
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1685868990
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_181
timestamp 1685868990
transform 1 0 17756 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1685868990
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1685868990
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_197
timestamp 1685868990
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_212
timestamp 1685868990
transform 1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1685868990
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1685868990
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_232
timestamp 1685868990
transform 1 0 22448 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_236
timestamp 1685868990
transform 1 0 22816 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1685868990
transform 1 0 23460 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_250
timestamp 1685868990
transform 1 0 24104 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_253
timestamp 1685868990
transform 1 0 24380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1685868990
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_269
timestamp 1685868990
transform 1 0 25852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1685868990
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1685868990
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1685868990
transform 1 0 27416 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1685868990
transform 1 0 28060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_300
timestamp 1685868990
transform 1 0 28704 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_309
timestamp 1685868990
transform 1 0 29532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_314
timestamp 1685868990
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_321
timestamp 1685868990
transform 1 0 30636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1685868990
transform 1 0 31740 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_337
timestamp 1685868990
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1685868990
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1685868990
transform -1 0 32476 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1685868990
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1685868990
transform -1 0 32476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1685868990
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1685868990
transform -1 0 32476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1685868990
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1685868990
transform -1 0 32476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1685868990
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1685868990
transform -1 0 32476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1685868990
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1685868990
transform -1 0 32476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1685868990
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1685868990
transform -1 0 32476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1685868990
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1685868990
transform -1 0 32476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1685868990
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1685868990
transform -1 0 32476 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1685868990
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1685868990
transform -1 0 32476 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1685868990
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1685868990
transform -1 0 32476 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1685868990
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1685868990
transform -1 0 32476 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1685868990
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1685868990
transform -1 0 32476 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1685868990
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1685868990
transform -1 0 32476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1685868990
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1685868990
transform -1 0 32476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1685868990
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1685868990
transform -1 0 32476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1685868990
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1685868990
transform -1 0 32476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1685868990
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1685868990
transform -1 0 32476 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1685868990
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1685868990
transform -1 0 32476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1685868990
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1685868990
transform -1 0 32476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1685868990
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1685868990
transform -1 0 32476 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1685868990
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1685868990
transform -1 0 32476 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1685868990
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1685868990
transform -1 0 32476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1685868990
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1685868990
transform -1 0 32476 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1685868990
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1685868990
transform -1 0 32476 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1685868990
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1685868990
transform -1 0 32476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1685868990
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1685868990
transform -1 0 32476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1685868990
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1685868990
transform -1 0 32476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1685868990
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1685868990
transform -1 0 32476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1685868990
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1685868990
transform -1 0 32476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1685868990
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1685868990
transform -1 0 32476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1685868990
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1685868990
transform -1 0 32476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1685868990
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1685868990
transform -1 0 32476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1685868990
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1685868990
transform -1 0 32476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1685868990
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1685868990
transform -1 0 32476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1685868990
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1685868990
transform -1 0 32476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1685868990
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1685868990
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1685868990
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1685868990
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1685868990
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1685868990
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1685868990
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1685868990
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1685868990
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1685868990
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1685868990
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1685868990
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1685868990
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1685868990
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1685868990
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1685868990
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1685868990
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1685868990
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1685868990
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1685868990
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1685868990
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1685868990
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1685868990
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1685868990
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1685868990
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1685868990
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1685868990
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1685868990
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1685868990
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1685868990
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1685868990
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1685868990
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1685868990
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1685868990
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1685868990
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1685868990
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1685868990
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1685868990
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1685868990
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1685868990
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1685868990
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1685868990
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1685868990
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1685868990
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1685868990
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1685868990
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1685868990
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1685868990
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1685868990
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1685868990
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1685868990
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1685868990
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1685868990
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1685868990
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1685868990
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1685868990
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1685868990
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1685868990
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1685868990
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1685868990
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1685868990
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1685868990
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1685868990
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1685868990
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1685868990
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1685868990
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1685868990
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1685868990
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1685868990
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1685868990
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1685868990
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1685868990
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1685868990
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1685868990
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1685868990
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1685868990
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1685868990
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1685868990
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1685868990
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1685868990
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1685868990
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1685868990
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1685868990
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1685868990
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1685868990
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1685868990
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1685868990
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1685868990
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1685868990
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1685868990
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1685868990
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1685868990
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1685868990
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1685868990
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1685868990
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1685868990
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1685868990
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1685868990
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1685868990
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1685868990
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1685868990
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1685868990
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1685868990
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1685868990
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1685868990
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1685868990
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1685868990
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1685868990
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1685868990
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1685868990
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1685868990
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1685868990
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1685868990
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1685868990
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1685868990
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1685868990
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1685868990
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1685868990
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1685868990
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1685868990
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1685868990
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1685868990
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1685868990
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1685868990
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1685868990
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1685868990
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1685868990
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1685868990
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1685868990
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1685868990
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1685868990
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1685868990
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1685868990
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1685868990
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1685868990
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1685868990
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1685868990
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1685868990
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1685868990
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1685868990
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1685868990
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1685868990
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1685868990
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1685868990
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1685868990
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1685868990
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1685868990
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1685868990
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1685868990
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1685868990
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1685868990
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1685868990
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1685868990
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1685868990
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1685868990
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1685868990
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1685868990
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1685868990
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1685868990
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1685868990
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1685868990
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1685868990
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1685868990
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1685868990
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1685868990
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1685868990
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1685868990
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1685868990
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1685868990
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1685868990
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1685868990
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1685868990
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1685868990
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1685868990
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1685868990
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1685868990
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1685868990
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1685868990
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1685868990
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1685868990
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1685868990
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1685868990
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1685868990
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1685868990
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1685868990
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1685868990
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1685868990
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1685868990
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1685868990
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1685868990
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1685868990
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1685868990
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1685868990
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1685868990
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1685868990
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1685868990
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1685868990
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1685868990
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1685868990
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1685868990
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1685868990
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1685868990
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1685868990
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1685868990
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1685868990
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1685868990
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1685868990
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1685868990
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1685868990
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1685868990
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1685868990
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1685868990
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1685868990
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1685868990
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1685868990
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1685868990
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1685868990
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1685868990
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1685868990
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1685868990
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1685868990
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1685868990
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1685868990
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1685868990
transform 1 0 24288 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1685868990
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1685868990
transform 1 0 29440 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1685868990
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_2  _31_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 23092 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _32_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 23368 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _33_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 23460 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _34_
timestamp 1685868990
transform -1 0 23276 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _35_
timestamp 1685868990
transform -1 0 25116 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _36_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 24288 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _37_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _38_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 21528 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_4  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 20608 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _40_
timestamp 1685868990
transform -1 0 22264 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 24656 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _42_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 23644 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _43_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 19872 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_4  _44_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 21988 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _45_
timestamp 1685868990
transform 1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _46_
timestamp 1685868990
transform -1 0 22356 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_2  _47_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 25208 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _48_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 22724 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _49_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 10948 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  _50_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 23736 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _51_
timestamp 1685868990
transform -1 0 21896 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _52_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 18860 0 -1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__o21a_1  _53_
timestamp 1685868990
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _54_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 18492 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _55_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 17480 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _56_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 24104 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _57_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 20976 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _58_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _59_
timestamp 1685868990
transform -1 0 22448 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _60_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 25576 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _61_
timestamp 1685868990
transform -1 0 17204 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__or2b_2  _62_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 24472 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _63_
timestamp 1685868990
transform -1 0 18308 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _64_
timestamp 1685868990
transform 1 0 11776 0 -1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_2  _65_
timestamp 1685868990
transform -1 0 11684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _66_
timestamp 1685868990
transform 1 0 6532 0 -1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _67_
timestamp 1685868990
transform -1 0 25944 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _68_
timestamp 1685868990
transform 1 0 20148 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1685868990
transform 1 0 20700 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 30360 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1685868990
transform 1 0 29716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1685868990
transform 1 0 28796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1685868990
transform 1 0 28428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1685868990
transform 1 0 27784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1685868990
transform 1 0 27140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1685868990
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1685868990
transform -1 0 25484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1685868990
transform 1 0 25576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1685868990
transform 1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1685868990
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1685868990
transform 1 0 23828 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1685868990
transform -1 0 20976 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1685868990
transform -1 0 18952 0 -1 20672
box -38 -48 314 592
use power_gate  power_gate_0 sky130_power_gate
timestamp 1685868990
transform 1 0 2670 0 1 -1530
box -1428 -1134 11168 908
use sky130_fd_sc_hd__conb_1  tt_um_power_test_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform -1 0 6992 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_16
timestamp 1685868990
transform 1 0 5796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_17
timestamp 1685868990
transform -1 0 5428 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_18
timestamp 1685868990
transform -1 0 4784 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_19
timestamp 1685868990
transform 1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_20
timestamp 1685868990
transform 1 0 2576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_21
timestamp 1685868990
transform 1 0 1932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_22
timestamp 1685868990
transform -1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_23
timestamp 1685868990
transform -1 0 13064 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_24
timestamp 1685868990
transform -1 0 12144 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_25
timestamp 1685868990
transform 1 0 10580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_26
timestamp 1685868990
transform 1 0 9936 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_27
timestamp 1685868990
transform 1 0 9292 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_28
timestamp 1685868990
transform -1 0 9200 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_29
timestamp 1685868990
transform -1 0 8464 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  tt_um_power_test_30
timestamp 1685868990
transform -1 0 7728 0 1 19584
box -38 -48 314 592
<< labels >>
flabel metal4 s 31710 21560 31770 21760 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 32446 21560 32506 21760 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30974 21560 31034 21760 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30238 21560 30298 21760 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 29502 21560 29562 21760 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 28766 21560 28826 21760 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 28030 21560 28090 21760 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 27294 21560 27354 21760 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 26558 21560 26618 21760 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 25822 21560 25882 21760 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 25086 21560 25146 21760 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 24350 21560 24410 21760 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 23614 21560 23674 21760 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22878 21560 22938 21760 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 22142 21560 22202 21760 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21406 21560 21466 21760 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20670 21560 20730 21760 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 21560 19994 21760 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19198 21560 19258 21760 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 6686 21560 6746 21760 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal tristate
flabel metal4 s 5950 21560 6010 21760 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal tristate
flabel metal4 s 5214 21560 5274 21760 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal tristate
flabel metal4 s 4478 21560 4538 21760 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal tristate
flabel metal4 s 3742 21560 3802 21760 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal tristate
flabel metal4 s 3006 21560 3066 21760 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal tristate
flabel metal4 s 2270 21560 2330 21760 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal tristate
flabel metal4 s 1534 21560 1594 21760 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal tristate
flabel metal4 s 12574 21560 12634 21760 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal tristate
flabel metal4 s 11838 21560 11898 21760 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal tristate
flabel metal4 s 11102 21560 11162 21760 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal tristate
flabel metal4 s 10366 21560 10426 21760 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal tristate
flabel metal4 s 9630 21560 9690 21760 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal tristate
flabel metal4 s 8894 21560 8954 21760 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal tristate
flabel metal4 s 8158 21560 8218 21760 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal tristate
flabel metal4 s 7422 21560 7482 21760 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal tristate
flabel metal4 s 18462 21560 18522 21760 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal tristate
flabel metal4 s 17726 21560 17786 21760 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal tristate
flabel metal4 s 16990 21560 17050 21760 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal tristate
flabel metal4 s 16254 21560 16314 21760 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal tristate
flabel metal4 s 15518 21560 15578 21760 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal tristate
flabel metal4 s 14782 21560 14842 21760 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal tristate
flabel metal4 s 14046 21560 14106 21760 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal tristate
flabel metal4 s 13310 21560 13370 21760 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal tristate
flabel metal4 s 8786 1040 9106 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 16628 1040 16948 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 24470 1040 24790 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
flabel metal4 s 32312 1040 32632 20720 0 FreeSans 1920 90 0 0 vssd1
port 44 nsew ground bidirectional
rlabel metal1 16790 20128 16790 20128 0 vccd1
rlabel via1 16868 20672 16868 20672 0 vssd1
rlabel metal2 11454 19652 11454 19652 0 _00_
rlabel metal1 18078 20468 18078 20468 0 _01_
rlabel metal1 17618 19822 17618 19822 0 _02_
rlabel metal1 18906 20366 18906 20366 0 _03_
rlabel metal1 22034 12172 22034 12172 0 _04_
rlabel metal1 21804 12410 21804 12410 0 _05_
rlabel metal1 22908 12274 22908 12274 0 _06_
rlabel metal1 21298 12410 21298 12410 0 _07_
rlabel metal1 19872 20298 19872 20298 0 _08_
rlabel metal2 18078 20298 18078 20298 0 _09_
rlabel metal1 23414 17204 23414 17204 0 _10_
rlabel metal2 22402 18802 22402 18802 0 _11_
rlabel metal1 19504 19754 19504 19754 0 _12_
rlabel metal2 18262 20706 18262 20706 0 _13_
rlabel metal1 21758 19448 21758 19448 0 _14_
rlabel metal1 24426 18666 24426 18666 0 _15_
rlabel metal2 10258 19822 10258 19822 0 _16_
rlabel metal1 11638 19856 11638 19856 0 _17_
rlabel metal2 21850 19669 21850 19669 0 _18_
rlabel metal1 18722 19312 18722 19312 0 _19_
rlabel metal1 17848 16218 17848 16218 0 _20_
rlabel metal1 18446 19754 18446 19754 0 _21_
rlabel metal1 23966 19278 23966 19278 0 _22_
rlabel metal1 16974 19890 16974 19890 0 _23_
rlabel metal1 16514 18700 16514 18700 0 _24_
rlabel metal2 17066 18530 17066 18530 0 _25_
rlabel metal2 12466 16524 12466 16524 0 _26_
rlabel metal1 15548 20434 15548 20434 0 _27_
rlabel metal2 7590 20196 7590 20196 0 _28_
rlabel metal2 25530 14212 25530 14212 0 _29_
rlabel metal1 20516 14586 20516 14586 0 _30_
rlabel metal1 28152 13974 28152 13974 0 net1
rlabel metal2 23414 20196 23414 20196 0 net10
rlabel metal2 22770 19108 22770 19108 0 net11
rlabel metal1 23782 17646 23782 17646 0 net12
rlabel metal1 20378 19346 20378 19346 0 net13
rlabel metal2 18906 20128 18906 20128 0 net14
rlabel via2 6762 20043 6762 20043 0 net15
rlabel via2 6026 20451 6026 20451 0 net16
rlabel metal2 5198 20655 5198 20655 0 net17
rlabel via2 4554 20451 4554 20451 0 net18
rlabel via2 3450 20451 3450 20451 0 net19
rlabel metal1 24794 16524 24794 16524 0 net2
rlabel via2 2806 20451 2806 20451 0 net20
rlabel via2 2162 20451 2162 20451 0 net21
rlabel via2 1610 20043 1610 20043 0 net22
rlabel metal1 12742 20026 12742 20026 0 net23
rlabel metal2 11914 20349 11914 20349 0 net24
rlabel metal1 10948 20026 10948 20026 0 net25
rlabel via2 10166 20043 10166 20043 0 net26
rlabel metal1 9614 20026 9614 20026 0 net27
rlabel metal1 9062 19278 9062 19278 0 net28
rlabel via2 8234 20043 8234 20043 0 net29
rlabel metal1 23414 20434 23414 20434 0 net3
rlabel via2 7498 20043 7498 20043 0 net30
rlabel metal2 19826 20298 19826 20298 0 net4
rlabel metal1 23506 17680 23506 17680 0 net5
rlabel metal1 20746 19414 20746 19414 0 net6
rlabel metal1 23414 19890 23414 19890 0 net7
rlabel metal1 25576 13974 25576 13974 0 net8
rlabel metal1 24610 16592 24610 16592 0 net9
rlabel metal4 30268 21525 30268 21525 0 ui_in[0]
rlabel metal4 29532 21321 29532 21321 0 ui_in[1]
rlabel metal4 28796 21525 28796 21525 0 ui_in[2]
rlabel metal4 28060 21321 28060 21321 0 ui_in[3]
rlabel metal4 27324 21525 27324 21525 0 ui_in[4]
rlabel metal4 26588 21321 26588 21321 0 ui_in[5]
rlabel metal4 25852 21525 25852 21525 0 ui_in[6]
rlabel metal4 24380 21525 24380 21525 0 uio_in[0]
rlabel metal4 23644 21525 23644 21525 0 uio_in[1]
rlabel metal4 22908 21049 22908 21049 0 uio_in[2]
rlabel metal4 22172 21525 22172 21525 0 uio_in[3]
rlabel metal4 21436 21525 21436 21525 0 uio_in[4]
rlabel metal4 20700 21253 20700 21253 0 uio_in[5]
rlabel metal4 19964 21525 19964 21525 0 uio_in[6]
rlabel metal2 19274 21165 19274 21165 0 uo_out[0]
rlabel metal4 17756 21525 17756 21525 0 uo_out[1]
rlabel metal4 17020 21457 17020 21457 0 uo_out[2]
rlabel metal4 16284 21525 16284 21525 0 uo_out[3]
rlabel metal4 15548 21525 15548 21525 0 uo_out[4]
rlabel metal4 14812 21525 14812 21525 0 uo_out[5]
rlabel metal1 8510 20536 8510 20536 0 uo_out[6]
rlabel metal4 13340 21525 13340 21525 0 uo_out[7]
flabel metal4 -54 -330 590 20568 0 FreeSans 1600 0 0 0 vccd1
port 45 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 33580 21760
<< end >>
