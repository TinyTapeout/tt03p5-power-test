VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_power_test
  CLASS BLOCK ;
  FOREIGN tt_um_power_test ;
  ORIGIN 0.000 0.000 ;
  SIZE 167.900 BY 108.800 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 107.800 158.850 108.800 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 162.230 107.800 162.530 108.800 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 107.800 155.170 108.800 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 107.260 151.490 108.800 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 105.220 147.810 108.800 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 107.260 144.130 108.800 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 105.220 140.450 108.800 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 107.260 136.770 108.800 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 105.220 133.090 108.800 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 107.260 129.410 108.800 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 107.800 125.730 108.800 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 107.260 122.050 108.800 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 107.260 118.370 108.800 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 102.500 114.690 108.800 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 107.260 111.010 108.800 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 107.260 107.330 108.800 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 104.540 103.650 108.800 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 107.260 99.970 108.800 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 107.800 96.290 108.800 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 100.460 33.730 108.800 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 102.500 30.050 108.800 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 104.540 26.370 108.800 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 102.500 22.690 108.800 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 102.500 19.010 108.800 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 102.500 15.330 108.800 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 102.500 11.650 108.800 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 100.460 7.970 108.800 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 101.820 63.170 108.800 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 107.260 59.490 108.800 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 107.260 55.810 108.800 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 100.460 52.130 108.800 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 107.260 48.450 108.800 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 107.260 44.770 108.800 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 100.460 41.090 108.800 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 100.460 37.410 108.800 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 107.260 92.610 108.800 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 107.260 88.930 108.800 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 106.580 85.250 108.800 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 107.260 81.570 108.800 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 107.260 77.890 108.800 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 107.260 74.210 108.800 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 106.580 70.530 108.800 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 107.260 66.850 108.800 ;
    END
  END uo_out[7]
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 43.930 5.200 45.530 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 83.140 5.200 84.740 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 122.350 5.200 123.950 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 161.560 5.200 163.160 103.600 ;
    END
  END vssd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2.000 -8.000 4.000 100.600 ;
    END
  END vccd1
  OBS
      LAYER nwell ;
        RECT 5.175 -7.535 66.005 2.645 ;
      LAYER pwell ;
        RECT 66.025 -7.500 68.125 2.600 ;
      LAYER li1 ;
        RECT 5.355 0.000 162.380 103.445 ;
        RECT 5.355 -7.180 5.525 0.000 ;
        RECT 5.925 -6.465 6.095 0.000 ;
        RECT 6.405 -6.465 6.575 0.000 ;
        RECT 6.885 -6.465 7.055 0.000 ;
        RECT 7.365 -6.465 7.535 0.000 ;
        RECT 7.845 -6.465 8.015 0.000 ;
        RECT 8.325 -6.465 8.495 0.000 ;
        RECT 8.805 -6.465 8.975 0.000 ;
        RECT 9.285 -6.465 9.455 0.000 ;
        RECT 9.765 -6.465 9.935 0.000 ;
        RECT 10.245 -6.465 10.415 0.000 ;
        RECT 10.725 -6.465 10.895 0.000 ;
        RECT 11.205 -6.465 11.375 0.000 ;
        RECT 11.685 -6.465 11.855 0.000 ;
        RECT 12.165 -6.465 12.335 0.000 ;
        RECT 12.645 -6.465 12.815 0.000 ;
        RECT 13.125 -6.465 13.295 0.000 ;
        RECT 13.605 -6.465 13.775 0.000 ;
        RECT 14.085 -6.465 14.255 0.000 ;
        RECT 14.565 -6.465 14.735 0.000 ;
        RECT 15.045 -6.465 15.215 0.000 ;
        RECT 15.525 -6.465 15.695 0.000 ;
        RECT 16.005 -6.465 16.175 0.000 ;
        RECT 16.485 -6.465 16.655 0.000 ;
        RECT 16.965 -6.465 17.135 0.000 ;
        RECT 17.445 -6.465 17.615 0.000 ;
        RECT 17.925 -6.465 18.095 0.000 ;
        RECT 18.405 -6.465 18.575 0.000 ;
        RECT 18.885 -6.465 19.055 0.000 ;
        RECT 19.365 -6.465 19.535 0.000 ;
        RECT 19.845 -6.465 20.015 0.000 ;
        RECT 20.325 -6.465 20.495 0.000 ;
        RECT 20.805 -6.465 20.975 0.000 ;
        RECT 21.285 -6.465 21.455 0.000 ;
        RECT 21.765 -6.465 21.935 0.000 ;
        RECT 22.245 -6.465 22.415 0.000 ;
        RECT 22.725 -6.465 22.895 0.000 ;
        RECT 23.205 -6.465 23.375 0.000 ;
        RECT 23.685 -6.465 23.855 0.000 ;
        RECT 24.165 -6.465 24.335 0.000 ;
        RECT 24.645 -6.465 24.815 0.000 ;
        RECT 25.125 -6.465 25.295 0.000 ;
        RECT 25.605 -6.465 25.775 0.000 ;
        RECT 26.085 -6.465 26.255 0.000 ;
        RECT 26.565 -6.465 26.735 0.000 ;
        RECT 27.045 -6.465 27.215 0.000 ;
        RECT 27.525 -6.465 27.695 0.000 ;
        RECT 28.005 -6.465 28.175 0.000 ;
        RECT 28.485 -6.465 28.655 0.000 ;
        RECT 28.965 -6.465 29.135 0.000 ;
        RECT 29.445 -6.465 29.615 0.000 ;
        RECT 29.925 -6.465 30.095 0.000 ;
        RECT 30.405 -6.465 30.575 0.000 ;
        RECT 30.885 -6.465 31.055 0.000 ;
        RECT 31.365 -6.465 31.535 0.000 ;
        RECT 31.845 -6.465 32.015 0.000 ;
        RECT 32.325 -6.465 32.495 0.000 ;
        RECT 32.805 -6.465 32.975 0.000 ;
        RECT 33.285 -6.465 33.455 0.000 ;
        RECT 33.765 -6.465 33.935 0.000 ;
        RECT 34.245 -6.465 34.415 0.000 ;
        RECT 34.715 -6.465 34.885 0.000 ;
        RECT 35.195 -6.465 35.365 0.000 ;
        RECT 35.675 -6.465 35.845 0.000 ;
        RECT 36.155 -6.465 36.325 0.000 ;
        RECT 36.635 -6.465 36.805 0.000 ;
        RECT 37.115 -6.465 37.285 0.000 ;
        RECT 37.595 -6.465 37.765 0.000 ;
        RECT 38.075 -6.465 38.245 0.000 ;
        RECT 38.555 -6.465 38.725 0.000 ;
        RECT 39.035 -6.465 39.205 0.000 ;
        RECT 39.515 -6.465 39.685 0.000 ;
        RECT 39.995 -6.465 40.165 0.000 ;
        RECT 40.475 -6.465 40.645 0.000 ;
        RECT 40.955 -6.465 41.125 0.000 ;
        RECT 41.435 -6.465 41.605 0.000 ;
        RECT 41.915 -6.465 42.085 0.000 ;
        RECT 42.395 -6.465 42.565 0.000 ;
        RECT 42.875 -6.465 43.045 0.000 ;
        RECT 43.355 -6.465 43.525 0.000 ;
        RECT 43.835 -6.465 44.005 0.000 ;
        RECT 44.315 -6.465 44.485 0.000 ;
        RECT 44.795 -6.465 44.965 0.000 ;
        RECT 45.275 -6.465 45.445 0.000 ;
        RECT 45.755 -6.465 45.925 0.000 ;
        RECT 46.235 -6.465 46.405 0.000 ;
        RECT 46.715 -6.465 46.885 0.000 ;
        RECT 47.195 -6.465 47.365 0.000 ;
        RECT 47.675 -6.465 47.845 0.000 ;
        RECT 48.155 -6.465 48.325 0.000 ;
        RECT 48.635 -6.465 48.805 0.000 ;
        RECT 49.115 -6.465 49.285 0.000 ;
        RECT 49.595 -6.465 49.765 0.000 ;
        RECT 50.075 -6.465 50.245 0.000 ;
        RECT 50.555 -6.465 50.725 0.000 ;
        RECT 51.035 -6.465 51.205 0.000 ;
        RECT 51.515 -6.465 51.685 0.000 ;
        RECT 51.995 -6.465 52.165 0.000 ;
        RECT 52.475 -6.465 52.645 0.000 ;
        RECT 52.955 -6.465 53.125 0.000 ;
        RECT 53.435 -6.465 53.605 0.000 ;
        RECT 53.915 -6.465 54.085 0.000 ;
        RECT 54.395 -6.465 54.565 0.000 ;
        RECT 54.875 -6.465 55.045 0.000 ;
        RECT 55.355 -6.465 55.525 0.000 ;
        RECT 55.835 -6.465 56.005 0.000 ;
        RECT 56.315 -6.465 56.485 0.000 ;
        RECT 56.795 -6.465 56.965 0.000 ;
        RECT 57.275 -6.465 57.445 0.000 ;
        RECT 57.755 -6.465 57.925 0.000 ;
        RECT 58.235 -6.465 58.405 0.000 ;
        RECT 58.715 -6.465 58.885 0.000 ;
        RECT 59.195 -6.465 59.365 0.000 ;
        RECT 59.675 -6.465 59.845 0.000 ;
        RECT 60.155 -6.465 60.325 0.000 ;
        RECT 60.635 -6.465 60.805 0.000 ;
        RECT 61.115 -6.465 61.285 0.000 ;
        RECT 61.595 -6.465 61.765 0.000 ;
        RECT 62.075 -6.465 62.245 0.000 ;
        RECT 62.555 -6.465 62.725 0.000 ;
        RECT 63.035 -6.465 63.205 0.000 ;
        RECT 63.515 -6.465 63.685 0.000 ;
        RECT 64.085 -6.465 64.815 0.000 ;
        RECT 65.085 -6.465 65.255 0.000 ;
        RECT 64.085 -6.470 64.780 -6.465 ;
        RECT 6.085 -6.855 6.415 -6.685 ;
        RECT 7.045 -6.855 7.375 -6.685 ;
        RECT 8.005 -6.855 8.335 -6.685 ;
        RECT 8.965 -6.855 9.295 -6.685 ;
        RECT 9.925 -6.855 10.255 -6.685 ;
        RECT 10.885 -6.855 11.215 -6.685 ;
        RECT 11.845 -6.855 12.175 -6.685 ;
        RECT 12.805 -6.855 13.135 -6.685 ;
        RECT 13.765 -6.855 14.095 -6.685 ;
        RECT 14.725 -6.855 15.055 -6.685 ;
        RECT 15.685 -6.855 16.015 -6.685 ;
        RECT 16.645 -6.855 16.975 -6.685 ;
        RECT 17.605 -6.855 17.935 -6.685 ;
        RECT 18.565 -6.855 18.895 -6.685 ;
        RECT 19.525 -6.855 19.855 -6.685 ;
        RECT 20.485 -6.855 20.815 -6.685 ;
        RECT 21.445 -6.855 21.775 -6.685 ;
        RECT 22.405 -6.855 22.735 -6.685 ;
        RECT 23.365 -6.855 23.695 -6.685 ;
        RECT 24.325 -6.855 24.655 -6.685 ;
        RECT 25.285 -6.855 25.615 -6.685 ;
        RECT 26.245 -6.855 26.575 -6.685 ;
        RECT 27.205 -6.855 27.535 -6.685 ;
        RECT 28.165 -6.855 28.495 -6.685 ;
        RECT 29.125 -6.855 29.455 -6.685 ;
        RECT 30.085 -6.855 30.415 -6.685 ;
        RECT 31.045 -6.855 31.375 -6.685 ;
        RECT 32.005 -6.855 32.335 -6.685 ;
        RECT 32.965 -6.855 33.295 -6.685 ;
        RECT 33.925 -6.855 34.255 -6.685 ;
        RECT 34.875 -6.855 35.205 -6.685 ;
        RECT 35.835 -6.855 36.165 -6.685 ;
        RECT 36.795 -6.855 37.125 -6.685 ;
        RECT 37.755 -6.855 38.085 -6.685 ;
        RECT 38.715 -6.855 39.045 -6.685 ;
        RECT 39.675 -6.855 40.005 -6.685 ;
        RECT 40.635 -6.855 40.965 -6.685 ;
        RECT 41.595 -6.855 41.925 -6.685 ;
        RECT 42.555 -6.855 42.885 -6.685 ;
        RECT 43.515 -6.855 43.845 -6.685 ;
        RECT 44.475 -6.855 44.805 -6.685 ;
        RECT 45.435 -6.855 45.765 -6.685 ;
        RECT 46.395 -6.855 46.725 -6.685 ;
        RECT 47.355 -6.855 47.685 -6.685 ;
        RECT 48.315 -6.855 48.645 -6.685 ;
        RECT 49.275 -6.855 49.605 -6.685 ;
        RECT 50.235 -6.855 50.565 -6.685 ;
        RECT 51.195 -6.855 51.525 -6.685 ;
        RECT 52.155 -6.855 52.485 -6.685 ;
        RECT 53.115 -6.855 53.445 -6.685 ;
        RECT 54.075 -6.855 54.405 -6.685 ;
        RECT 55.035 -6.855 55.365 -6.685 ;
        RECT 55.995 -6.855 56.325 -6.685 ;
        RECT 56.955 -6.855 57.285 -6.685 ;
        RECT 57.915 -6.855 58.245 -6.685 ;
        RECT 58.875 -6.855 59.205 -6.685 ;
        RECT 59.835 -6.855 60.165 -6.685 ;
        RECT 60.795 -6.855 61.125 -6.685 ;
        RECT 61.755 -6.855 62.085 -6.685 ;
        RECT 62.715 -6.855 63.045 -6.685 ;
        RECT 64.085 -7.180 64.255 -6.470 ;
        RECT 64.785 -6.895 65.165 -6.695 ;
        RECT 65.655 -7.180 65.825 0.000 ;
        RECT 5.355 -7.355 65.825 -7.180 ;
        RECT 66.205 -7.150 66.375 0.000 ;
        RECT 66.755 -6.470 66.925 0.000 ;
        RECT 67.225 -1.540 67.950 0.000 ;
        RECT 67.225 -6.460 67.945 -1.540 ;
        RECT 67.225 -6.470 67.395 -6.460 ;
        RECT 66.865 -6.810 67.295 -6.640 ;
        RECT 67.775 -7.150 67.945 -6.460 ;
        RECT 66.205 -7.320 67.945 -7.150 ;
        RECT 5.510 -7.360 65.670 -7.355 ;
      LAYER met1 ;
        RECT 5.450 0.000 164.600 106.580 ;
        RECT 5.810 -1.440 6.200 0.000 ;
        RECT 5.895 -6.445 6.125 -1.440 ;
        RECT 6.375 -3.440 6.605 0.000 ;
        RECT 6.770 -1.440 7.160 0.000 ;
        RECT 6.290 -6.440 6.680 -3.440 ;
        RECT 6.375 -6.445 6.605 -6.440 ;
        RECT 6.855 -6.445 7.085 -1.440 ;
        RECT 7.335 -3.440 7.565 0.000 ;
        RECT 7.730 -1.440 8.120 0.000 ;
        RECT 7.250 -6.440 7.640 -3.440 ;
        RECT 7.335 -6.445 7.565 -6.440 ;
        RECT 7.815 -6.445 8.045 -1.440 ;
        RECT 8.295 -3.440 8.525 0.000 ;
        RECT 8.690 -1.440 9.080 0.000 ;
        RECT 8.210 -6.440 8.600 -3.440 ;
        RECT 8.295 -6.445 8.525 -6.440 ;
        RECT 8.775 -6.445 9.005 -1.440 ;
        RECT 9.255 -3.440 9.485 0.000 ;
        RECT 9.650 -1.440 10.040 0.000 ;
        RECT 9.170 -6.440 9.560 -3.440 ;
        RECT 9.255 -6.445 9.485 -6.440 ;
        RECT 9.735 -6.445 9.965 -1.440 ;
        RECT 10.215 -3.440 10.445 0.000 ;
        RECT 10.610 -1.440 11.000 0.000 ;
        RECT 10.130 -6.440 10.520 -3.440 ;
        RECT 10.215 -6.445 10.445 -6.440 ;
        RECT 10.695 -6.445 10.925 -1.440 ;
        RECT 11.175 -3.440 11.405 0.000 ;
        RECT 11.570 -1.440 11.960 0.000 ;
        RECT 11.090 -6.440 11.480 -3.440 ;
        RECT 11.175 -6.445 11.405 -6.440 ;
        RECT 11.655 -6.445 11.885 -1.440 ;
        RECT 12.135 -3.440 12.365 0.000 ;
        RECT 12.530 -1.440 12.920 0.000 ;
        RECT 12.050 -6.440 12.440 -3.440 ;
        RECT 12.135 -6.445 12.365 -6.440 ;
        RECT 12.615 -6.445 12.845 -1.440 ;
        RECT 13.095 -3.440 13.325 0.000 ;
        RECT 13.490 -1.440 13.880 0.000 ;
        RECT 13.010 -6.440 13.400 -3.440 ;
        RECT 13.095 -6.445 13.325 -6.440 ;
        RECT 13.575 -6.445 13.805 -1.440 ;
        RECT 14.055 -3.440 14.285 0.000 ;
        RECT 14.450 -1.440 14.840 0.000 ;
        RECT 13.970 -6.440 14.360 -3.440 ;
        RECT 14.055 -6.445 14.285 -6.440 ;
        RECT 14.535 -6.445 14.765 -1.440 ;
        RECT 15.015 -3.440 15.245 0.000 ;
        RECT 15.410 -1.440 15.800 0.000 ;
        RECT 14.930 -6.440 15.320 -3.440 ;
        RECT 15.015 -6.445 15.245 -6.440 ;
        RECT 15.495 -6.445 15.725 -1.440 ;
        RECT 15.975 -3.440 16.205 0.000 ;
        RECT 16.370 -1.440 16.760 0.000 ;
        RECT 15.890 -6.440 16.280 -3.440 ;
        RECT 15.975 -6.445 16.205 -6.440 ;
        RECT 16.455 -6.445 16.685 -1.440 ;
        RECT 16.935 -3.440 17.165 0.000 ;
        RECT 17.330 -1.440 17.720 0.000 ;
        RECT 16.850 -6.440 17.240 -3.440 ;
        RECT 16.935 -6.445 17.165 -6.440 ;
        RECT 17.415 -6.445 17.645 -1.440 ;
        RECT 17.895 -3.440 18.125 0.000 ;
        RECT 18.290 -1.440 18.680 0.000 ;
        RECT 17.810 -6.440 18.200 -3.440 ;
        RECT 17.895 -6.445 18.125 -6.440 ;
        RECT 18.375 -6.445 18.605 -1.440 ;
        RECT 18.855 -3.440 19.085 0.000 ;
        RECT 19.250 -1.440 19.640 0.000 ;
        RECT 18.770 -6.440 19.160 -3.440 ;
        RECT 18.855 -6.445 19.085 -6.440 ;
        RECT 19.335 -6.445 19.565 -1.440 ;
        RECT 19.815 -3.440 20.045 0.000 ;
        RECT 20.210 -1.440 20.600 0.000 ;
        RECT 19.730 -6.440 20.120 -3.440 ;
        RECT 19.815 -6.445 20.045 -6.440 ;
        RECT 20.295 -6.445 20.525 -1.440 ;
        RECT 20.775 -3.440 21.005 0.000 ;
        RECT 21.170 -1.440 21.560 0.000 ;
        RECT 20.690 -6.440 21.080 -3.440 ;
        RECT 20.775 -6.445 21.005 -6.440 ;
        RECT 21.255 -6.445 21.485 -1.440 ;
        RECT 21.735 -3.440 21.965 0.000 ;
        RECT 22.130 -1.440 22.520 0.000 ;
        RECT 21.650 -6.440 22.040 -3.440 ;
        RECT 21.735 -6.445 21.965 -6.440 ;
        RECT 22.215 -6.445 22.445 -1.440 ;
        RECT 22.695 -3.440 22.925 0.000 ;
        RECT 23.090 -1.440 23.480 0.000 ;
        RECT 22.610 -6.440 23.000 -3.440 ;
        RECT 22.695 -6.445 22.925 -6.440 ;
        RECT 23.175 -6.445 23.405 -1.440 ;
        RECT 23.655 -3.440 23.885 0.000 ;
        RECT 24.050 -1.440 24.440 0.000 ;
        RECT 23.570 -6.440 23.960 -3.440 ;
        RECT 23.655 -6.445 23.885 -6.440 ;
        RECT 24.135 -6.445 24.365 -1.440 ;
        RECT 24.615 -3.440 24.845 0.000 ;
        RECT 25.010 -1.440 25.400 0.000 ;
        RECT 24.530 -6.440 24.920 -3.440 ;
        RECT 24.615 -6.445 24.845 -6.440 ;
        RECT 25.095 -6.445 25.325 -1.440 ;
        RECT 25.575 -3.440 25.805 0.000 ;
        RECT 25.970 -1.440 26.360 0.000 ;
        RECT 25.490 -6.440 25.880 -3.440 ;
        RECT 25.575 -6.445 25.805 -6.440 ;
        RECT 26.055 -6.445 26.285 -1.440 ;
        RECT 26.535 -3.440 26.765 0.000 ;
        RECT 26.930 -1.440 27.320 0.000 ;
        RECT 26.450 -6.440 26.840 -3.440 ;
        RECT 26.535 -6.445 26.765 -6.440 ;
        RECT 27.015 -6.445 27.245 -1.440 ;
        RECT 27.495 -3.440 27.725 0.000 ;
        RECT 27.890 -1.440 28.280 0.000 ;
        RECT 27.410 -6.440 27.800 -3.440 ;
        RECT 27.495 -6.445 27.725 -6.440 ;
        RECT 27.975 -6.445 28.205 -1.440 ;
        RECT 28.455 -3.440 28.685 0.000 ;
        RECT 28.850 -1.440 29.240 0.000 ;
        RECT 28.370 -6.440 28.760 -3.440 ;
        RECT 28.455 -6.445 28.685 -6.440 ;
        RECT 28.935 -6.445 29.165 -1.440 ;
        RECT 29.415 -3.440 29.645 0.000 ;
        RECT 29.810 -1.440 30.200 0.000 ;
        RECT 29.330 -6.440 29.720 -3.440 ;
        RECT 29.415 -6.445 29.645 -6.440 ;
        RECT 29.895 -6.445 30.125 -1.440 ;
        RECT 30.375 -3.440 30.605 0.000 ;
        RECT 30.770 -1.440 31.160 0.000 ;
        RECT 30.290 -6.440 30.680 -3.440 ;
        RECT 30.375 -6.445 30.605 -6.440 ;
        RECT 30.855 -6.445 31.085 -1.440 ;
        RECT 31.335 -3.440 31.565 0.000 ;
        RECT 31.730 -1.440 32.120 0.000 ;
        RECT 31.250 -6.440 31.640 -3.440 ;
        RECT 31.335 -6.445 31.565 -6.440 ;
        RECT 31.815 -6.445 32.045 -1.440 ;
        RECT 32.295 -3.440 32.525 0.000 ;
        RECT 32.690 -1.440 33.080 0.000 ;
        RECT 32.210 -6.440 32.600 -3.440 ;
        RECT 32.295 -6.445 32.525 -6.440 ;
        RECT 32.775 -6.445 33.005 -1.440 ;
        RECT 33.255 -3.440 33.485 0.000 ;
        RECT 33.650 -1.440 34.040 0.000 ;
        RECT 33.170 -6.440 33.560 -3.440 ;
        RECT 33.255 -6.445 33.485 -6.440 ;
        RECT 33.735 -6.445 33.965 -1.440 ;
        RECT 34.215 -3.440 34.445 0.000 ;
        RECT 34.610 -1.440 35.000 0.000 ;
        RECT 34.130 -6.440 34.520 -3.440 ;
        RECT 34.215 -6.445 34.445 -6.440 ;
        RECT 34.685 -6.445 34.915 -1.440 ;
        RECT 35.165 -3.440 35.395 0.000 ;
        RECT 35.570 -1.440 35.960 0.000 ;
        RECT 35.090 -6.440 35.480 -3.440 ;
        RECT 35.165 -6.445 35.395 -6.440 ;
        RECT 35.645 -6.445 35.875 -1.440 ;
        RECT 36.125 -3.440 36.355 0.000 ;
        RECT 36.530 -1.440 36.920 0.000 ;
        RECT 36.050 -6.440 36.440 -3.440 ;
        RECT 36.125 -6.445 36.355 -6.440 ;
        RECT 36.605 -6.445 36.835 -1.440 ;
        RECT 37.085 -3.440 37.315 0.000 ;
        RECT 37.490 -1.440 37.880 0.000 ;
        RECT 37.010 -6.440 37.400 -3.440 ;
        RECT 37.085 -6.445 37.315 -6.440 ;
        RECT 37.565 -6.445 37.795 -1.440 ;
        RECT 38.045 -3.440 38.275 0.000 ;
        RECT 38.450 -1.440 38.840 0.000 ;
        RECT 37.970 -6.440 38.360 -3.440 ;
        RECT 38.045 -6.445 38.275 -6.440 ;
        RECT 38.525 -6.445 38.755 -1.440 ;
        RECT 39.005 -3.440 39.235 0.000 ;
        RECT 39.410 -1.440 39.800 0.000 ;
        RECT 38.930 -6.440 39.320 -3.440 ;
        RECT 39.005 -6.445 39.235 -6.440 ;
        RECT 39.485 -6.445 39.715 -1.440 ;
        RECT 39.965 -3.440 40.195 0.000 ;
        RECT 40.370 -1.440 40.760 0.000 ;
        RECT 39.890 -6.440 40.280 -3.440 ;
        RECT 39.965 -6.445 40.195 -6.440 ;
        RECT 40.445 -6.445 40.675 -1.440 ;
        RECT 40.925 -3.440 41.155 0.000 ;
        RECT 41.330 -1.440 41.720 0.000 ;
        RECT 40.850 -6.440 41.240 -3.440 ;
        RECT 40.925 -6.445 41.155 -6.440 ;
        RECT 41.405 -6.445 41.635 -1.440 ;
        RECT 41.885 -3.440 42.115 0.000 ;
        RECT 42.290 -1.440 42.680 0.000 ;
        RECT 41.810 -6.440 42.200 -3.440 ;
        RECT 41.885 -6.445 42.115 -6.440 ;
        RECT 42.365 -6.445 42.595 -1.440 ;
        RECT 42.845 -3.440 43.075 0.000 ;
        RECT 43.250 -1.440 43.640 0.000 ;
        RECT 42.770 -6.440 43.160 -3.440 ;
        RECT 42.845 -6.445 43.075 -6.440 ;
        RECT 43.325 -6.445 43.555 -1.440 ;
        RECT 43.805 -3.440 44.035 0.000 ;
        RECT 44.210 -1.440 44.600 0.000 ;
        RECT 43.730 -6.440 44.120 -3.440 ;
        RECT 43.805 -6.445 44.035 -6.440 ;
        RECT 44.285 -6.445 44.515 -1.440 ;
        RECT 44.765 -3.440 44.995 0.000 ;
        RECT 45.170 -1.440 45.560 0.000 ;
        RECT 44.690 -6.440 45.080 -3.440 ;
        RECT 44.765 -6.445 44.995 -6.440 ;
        RECT 45.245 -6.445 45.475 -1.440 ;
        RECT 45.725 -3.440 45.955 0.000 ;
        RECT 46.130 -1.440 46.520 0.000 ;
        RECT 45.650 -6.440 46.040 -3.440 ;
        RECT 45.725 -6.445 45.955 -6.440 ;
        RECT 46.205 -6.445 46.435 -1.440 ;
        RECT 46.685 -3.440 46.915 0.000 ;
        RECT 47.090 -1.440 47.480 0.000 ;
        RECT 46.610 -6.440 47.000 -3.440 ;
        RECT 46.685 -6.445 46.915 -6.440 ;
        RECT 47.165 -6.445 47.395 -1.440 ;
        RECT 47.645 -3.440 47.875 0.000 ;
        RECT 48.050 -1.440 48.440 0.000 ;
        RECT 47.570 -6.440 47.960 -3.440 ;
        RECT 47.645 -6.445 47.875 -6.440 ;
        RECT 48.125 -6.445 48.355 -1.440 ;
        RECT 48.605 -3.440 48.835 0.000 ;
        RECT 49.010 -1.440 49.400 0.000 ;
        RECT 48.530 -6.440 48.920 -3.440 ;
        RECT 48.605 -6.445 48.835 -6.440 ;
        RECT 49.085 -6.445 49.315 -1.440 ;
        RECT 49.565 -3.440 49.795 0.000 ;
        RECT 49.970 -1.440 50.360 0.000 ;
        RECT 49.490 -6.440 49.880 -3.440 ;
        RECT 49.565 -6.445 49.795 -6.440 ;
        RECT 50.045 -6.445 50.275 -1.440 ;
        RECT 50.525 -3.440 50.755 0.000 ;
        RECT 50.930 -1.440 51.320 0.000 ;
        RECT 50.450 -6.440 50.840 -3.440 ;
        RECT 50.525 -6.445 50.755 -6.440 ;
        RECT 51.005 -6.445 51.235 -1.440 ;
        RECT 51.485 -3.440 51.715 0.000 ;
        RECT 51.890 -1.440 52.280 0.000 ;
        RECT 51.410 -6.440 51.800 -3.440 ;
        RECT 51.485 -6.445 51.715 -6.440 ;
        RECT 51.965 -6.445 52.195 -1.440 ;
        RECT 52.445 -3.440 52.675 0.000 ;
        RECT 52.850 -1.440 53.240 0.000 ;
        RECT 52.370 -6.440 52.760 -3.440 ;
        RECT 52.445 -6.445 52.675 -6.440 ;
        RECT 52.925 -6.445 53.155 -1.440 ;
        RECT 53.405 -3.440 53.635 0.000 ;
        RECT 53.810 -1.440 54.200 0.000 ;
        RECT 53.330 -6.440 53.720 -3.440 ;
        RECT 53.405 -6.445 53.635 -6.440 ;
        RECT 53.885 -6.445 54.115 -1.440 ;
        RECT 54.365 -3.440 54.595 0.000 ;
        RECT 54.770 -1.440 55.160 0.000 ;
        RECT 54.290 -6.440 54.680 -3.440 ;
        RECT 54.365 -6.445 54.595 -6.440 ;
        RECT 54.845 -6.445 55.075 -1.440 ;
        RECT 55.325 -3.450 55.555 0.000 ;
        RECT 55.730 -1.440 56.120 0.000 ;
        RECT 55.250 -6.450 55.640 -3.450 ;
        RECT 55.805 -6.445 56.035 -1.440 ;
        RECT 56.285 -3.450 56.515 0.000 ;
        RECT 56.690 -1.440 57.080 0.000 ;
        RECT 56.210 -6.450 56.600 -3.450 ;
        RECT 56.765 -6.445 56.995 -1.440 ;
        RECT 57.245 -3.450 57.475 0.000 ;
        RECT 57.650 -1.440 58.040 0.000 ;
        RECT 57.170 -6.450 57.560 -3.450 ;
        RECT 57.725 -6.445 57.955 -1.440 ;
        RECT 58.205 -3.450 58.435 0.000 ;
        RECT 58.610 -1.440 59.000 0.000 ;
        RECT 58.130 -6.450 58.520 -3.450 ;
        RECT 58.685 -6.445 58.915 -1.440 ;
        RECT 59.165 -3.450 59.395 0.000 ;
        RECT 59.570 -1.440 59.960 0.000 ;
        RECT 59.090 -6.450 59.480 -3.450 ;
        RECT 59.645 -6.445 59.875 -1.440 ;
        RECT 60.125 -3.450 60.355 0.000 ;
        RECT 60.530 -1.440 60.920 0.000 ;
        RECT 60.050 -6.450 60.440 -3.450 ;
        RECT 60.605 -6.445 60.835 -1.440 ;
        RECT 61.085 -3.450 61.315 0.000 ;
        RECT 61.490 -1.440 61.880 0.000 ;
        RECT 61.010 -6.450 61.400 -3.450 ;
        RECT 61.565 -6.445 61.795 -1.440 ;
        RECT 62.045 -3.450 62.275 0.000 ;
        RECT 62.450 -1.440 62.840 0.000 ;
        RECT 61.970 -6.450 62.360 -3.450 ;
        RECT 62.525 -6.445 62.755 -1.440 ;
        RECT 63.005 -3.450 63.235 0.000 ;
        RECT 63.410 -1.440 63.800 0.000 ;
        RECT 62.930 -6.450 63.320 -3.450 ;
        RECT 63.485 -6.445 63.715 -1.440 ;
        RECT 64.010 -1.860 64.250 0.000 ;
        RECT 63.960 -3.100 64.470 -1.860 ;
        RECT 64.010 -6.650 64.250 -3.100 ;
        RECT 64.615 -3.390 64.845 0.000 ;
        RECT 64.490 -6.450 64.900 -3.390 ;
        RECT 65.055 -6.445 66.955 0.000 ;
        RECT 65.180 -6.450 66.955 -6.445 ;
        RECT 67.195 -1.600 68.000 0.000 ;
        RECT 67.195 -6.450 67.425 -1.600 ;
        RECT 6.100 -6.890 64.250 -6.650 ;
        RECT 64.720 -6.760 67.285 -6.610 ;
        RECT 64.725 -6.840 67.285 -6.760 ;
        RECT 64.725 -6.880 67.220 -6.840 ;
        RECT 64.725 -6.915 65.185 -6.880 ;
        RECT 5.460 -7.070 64.540 -7.050 ;
        RECT 5.460 -7.150 65.720 -7.070 ;
        RECT 5.450 -7.390 65.730 -7.150 ;
      LAYER met2 ;
        RECT 5.510 0.000 164.590 107.285 ;
        RECT 5.860 -1.540 63.750 0.000 ;
        RECT 67.630 -1.590 67.950 0.000 ;
        RECT 64.010 -3.160 65.890 -1.810 ;
        RECT 6.330 -6.540 63.270 -3.350 ;
        RECT 64.540 -7.000 64.850 -3.340 ;
        RECT 5.510 -7.410 65.670 -7.000 ;
      LAYER met3 ;
        RECT 5.160 0.000 164.670 107.265 ;
        RECT 5.160 -1.540 66.030 0.000 ;
        RECT 66.440 -1.540 68.130 0.000 ;
        RECT 5.250 -1.640 66.000 -1.540 ;
        RECT 66.480 -1.610 68.020 -1.540 ;
        RECT 5.170 -3.375 6.330 -3.370 ;
        RECT 5.170 -3.400 63.320 -3.375 ;
        RECT 5.170 -7.540 68.140 -3.400 ;
        RECT 5.330 -8.000 67.870 -7.540 ;
      LAYER met4 ;
        RECT 4.000 101.000 7.270 108.470 ;
        RECT 4.400 100.060 7.270 101.000 ;
        RECT 8.370 102.100 10.950 108.470 ;
        RECT 12.050 102.100 14.630 108.470 ;
        RECT 15.730 102.100 18.310 108.470 ;
        RECT 19.410 102.100 21.990 108.470 ;
        RECT 23.090 104.140 25.670 108.470 ;
        RECT 26.770 104.140 29.350 108.470 ;
        RECT 23.090 102.100 29.350 104.140 ;
        RECT 30.450 102.100 33.030 108.470 ;
        RECT 8.370 100.060 33.030 102.100 ;
        RECT 34.130 100.060 36.710 108.470 ;
        RECT 37.810 100.060 40.390 108.470 ;
        RECT 41.490 106.860 44.070 108.470 ;
        RECT 45.170 106.860 47.750 108.470 ;
        RECT 48.850 106.860 51.430 108.470 ;
        RECT 41.490 104.000 51.430 106.860 ;
        RECT 41.490 100.060 43.530 104.000 ;
        RECT 4.400 4.800 43.530 100.060 ;
        RECT 45.930 100.060 51.430 104.000 ;
        RECT 52.530 106.860 55.110 108.470 ;
        RECT 56.210 106.860 58.790 108.470 ;
        RECT 59.890 106.860 62.470 108.470 ;
        RECT 52.530 101.420 62.470 106.860 ;
        RECT 63.570 106.860 66.150 108.470 ;
        RECT 67.250 106.860 69.830 108.470 ;
        RECT 63.570 106.180 69.830 106.860 ;
        RECT 70.930 106.860 73.510 108.470 ;
        RECT 74.610 106.860 77.190 108.470 ;
        RECT 78.290 106.860 80.870 108.470 ;
        RECT 81.970 106.860 84.550 108.470 ;
        RECT 70.930 106.180 84.550 106.860 ;
        RECT 85.650 106.860 88.230 108.470 ;
        RECT 89.330 106.860 91.910 108.470 ;
        RECT 93.010 107.400 95.590 108.470 ;
        RECT 96.690 107.400 99.270 108.470 ;
        RECT 93.010 106.860 99.270 107.400 ;
        RECT 100.370 106.860 102.950 108.470 ;
        RECT 85.650 106.180 102.950 106.860 ;
        RECT 63.570 104.140 102.950 106.180 ;
        RECT 104.050 106.860 106.630 108.470 ;
        RECT 107.730 106.860 110.310 108.470 ;
        RECT 111.410 106.860 113.990 108.470 ;
        RECT 104.050 104.140 113.990 106.860 ;
        RECT 63.570 104.000 113.990 104.140 ;
        RECT 63.570 101.420 82.740 104.000 ;
        RECT 52.530 100.060 82.740 101.420 ;
        RECT 45.930 4.800 82.740 100.060 ;
        RECT 85.140 102.100 113.990 104.000 ;
        RECT 115.090 106.860 117.670 108.470 ;
        RECT 118.770 106.860 121.350 108.470 ;
        RECT 122.450 107.400 125.030 108.470 ;
        RECT 126.130 107.400 128.710 108.470 ;
        RECT 122.450 106.860 128.710 107.400 ;
        RECT 129.810 106.860 132.390 108.470 ;
        RECT 115.090 104.820 132.390 106.860 ;
        RECT 133.490 106.860 136.070 108.470 ;
        RECT 137.170 106.860 139.750 108.470 ;
        RECT 133.490 104.820 139.750 106.860 ;
        RECT 140.850 106.860 143.430 108.470 ;
        RECT 144.530 106.860 147.110 108.470 ;
        RECT 140.850 104.820 147.110 106.860 ;
        RECT 148.210 106.860 150.790 108.470 ;
        RECT 151.890 107.400 154.470 108.470 ;
        RECT 155.570 107.400 158.150 108.470 ;
        RECT 159.250 107.400 161.830 108.470 ;
        RECT 162.930 107.400 164.670 108.470 ;
        RECT 151.890 106.860 164.670 107.400 ;
        RECT 148.210 104.820 164.670 106.860 ;
        RECT 115.090 104.000 164.670 104.820 ;
        RECT 115.090 102.100 121.950 104.000 ;
        RECT 85.140 4.800 121.950 102.100 ;
        RECT 124.350 4.800 161.160 104.000 ;
        RECT 163.560 4.800 164.670 104.000 ;
        RECT 4.400 0.000 164.670 4.800 ;
        RECT 4.800 -1.640 66.000 0.000 ;
        RECT 66.480 -1.610 163.140 0.000 ;
        RECT 4.000 -8.000 67.870 -3.760 ;
  END
END tt_um_power_test
END LIBRARY

